module challenge ( clk, n_rst, en, next_byte, win, state );
  input [6:0] next_byte;
  input clk, n_rst, en;
  output win;
  output state;
  wire   n1234, n1236, n1238, n1240, n1242, n1244, n1246, n1248, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
         n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
         n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
         n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
         n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
         n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
         n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
         n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
         n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
         n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
         n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
         n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
         n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
         n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
         n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
         n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
         n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
         n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
         n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
         n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
         n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
         n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
         n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
         n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
         n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
         n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
         n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
         n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
         n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
         n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
         n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
         n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
         n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831,
         n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
         n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
         n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
         n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
         n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
         n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
         n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
         n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
         n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
         n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931,
         n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
         n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
         n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
         n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971,
         n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
         n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
         n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
         n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011,
         n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021,
         n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
         n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
         n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
         n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
         n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
         n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
         n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
         n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
         n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
         n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
         n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
         n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
         n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
         n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
         n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
         n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
         n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
         n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
         n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
         n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
         n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
         n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
         n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
         n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
         n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
         n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481;
  wire   [7:0] state;
  

  DFFSR \state_reg[0]  ( .D(n1248), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        state[0]) );
  DFFSR \state_reg[1]  ( .D(n1246), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        state[1]) );
  DFFSR \state_reg[3]  ( .D(n1244), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        state[3]) );
  DFFSR \state_reg[7]  ( .D(n1242), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        state[7]) );
  DFFSR \state_reg[6]  ( .D(n1240), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        state[6]) );
  DFFSR \state_reg[5]  ( .D(n1238), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        state[5]) );
  DFFSR \state_reg[4]  ( .D(n1236), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        state[4]) );
  DFFSR \state_reg[2]  ( .D(n1234), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        state[2]) );
  BUFX2 U1252 ( .A(n2062), .Y(n1250) );
  AND2X2 U1253 ( .A(n1633), .B(n1250), .Y(n1963) );
  INVX2 U1254 ( .A(n2185), .Y(n1251) );
  INVX2 U1255 ( .A(n1254), .Y(n1678) );
  INVX2 U1256 ( .A(n2116), .Y(n1252) );
  AND2X2 U1257 ( .A(n2072), .B(n1252), .Y(n2355) );
  AND2X2 U1258 ( .A(n1922), .B(n1252), .Y(n1930) );
  INVX2 U1259 ( .A(n1451), .Y(n1414) );
  INVX2 U1260 ( .A(n1637), .Y(n1633) );
  INVX2 U1261 ( .A(n2406), .Y(n1601) );
  INVX2 U1262 ( .A(n2440), .Y(n1986) );
  INVX2 U1263 ( .A(n1800), .Y(n1982) );
  NOR2X1 U1264 ( .A(n1253), .B(n1254), .Y(win) );
  OR2X1 U1265 ( .A(n1255), .B(n1256), .Y(n1248) );
  MUX2X1 U1266 ( .B(n1257), .A(n1258), .S(n1259), .Y(n1256) );
  OAI21X1 U1267 ( .A(n1260), .B(n1261), .C(n1262), .Y(n1257) );
  NOR2X1 U1268 ( .A(n1263), .B(n1264), .Y(n1262) );
  AOI21X1 U1269 ( .A(n1265), .B(n1266), .C(n1267), .Y(n1261) );
  OAI21X1 U1270 ( .A(n1268), .B(n1269), .C(n1270), .Y(n1265) );
  OAI21X1 U1271 ( .A(n1271), .B(n1272), .C(n1273), .Y(n1269) );
  NOR2X1 U1272 ( .A(n1274), .B(n1275), .Y(n1271) );
  OAI21X1 U1273 ( .A(n1276), .B(n1277), .C(n1278), .Y(n1275) );
  OAI21X1 U1274 ( .A(n1279), .B(n1280), .C(n1281), .Y(n1277) );
  AOI21X1 U1275 ( .A(n1282), .B(n1283), .C(n1284), .Y(n1279) );
  OAI21X1 U1276 ( .A(n1285), .B(n1286), .C(n1287), .Y(n1284) );
  NAND3X1 U1277 ( .A(n1288), .B(n1289), .C(n1290), .Y(n1282) );
  OAI21X1 U1278 ( .A(n1291), .B(n1292), .C(n1293), .Y(n1290) );
  INVX1 U1279 ( .A(n1294), .Y(n1291) );
  OAI21X1 U1280 ( .A(n1295), .B(n1296), .C(n1297), .Y(n1294) );
  AND2X1 U1281 ( .A(n1298), .B(n1299), .Y(n1297) );
  OAI21X1 U1282 ( .A(n1300), .B(n1301), .C(n1302), .Y(n1296) );
  OAI21X1 U1283 ( .A(n1303), .B(n1304), .C(n1305), .Y(n1301) );
  AND2X1 U1284 ( .A(n1306), .B(n1307), .Y(n1304) );
  OAI21X1 U1285 ( .A(n1308), .B(n1309), .C(n1310), .Y(n1307) );
  OAI21X1 U1286 ( .A(n1311), .B(n1312), .C(n1313), .Y(n1309) );
  NAND2X1 U1287 ( .A(n1314), .B(n1315), .Y(n1312) );
  AOI21X1 U1288 ( .A(n1316), .B(n1317), .C(n1318), .Y(n1311) );
  OAI21X1 U1289 ( .A(n1319), .B(n1320), .C(n1321), .Y(n1316) );
  AND2X1 U1290 ( .A(n1322), .B(n1323), .Y(n1321) );
  NAND2X1 U1291 ( .A(n1324), .B(n1325), .Y(n1320) );
  OAI21X1 U1292 ( .A(n1326), .B(n1327), .C(n1328), .Y(n1324) );
  AOI21X1 U1293 ( .A(n1329), .B(n1330), .C(n1331), .Y(n1327) );
  NAND2X1 U1294 ( .A(n1332), .B(n1333), .Y(n1331) );
  OAI21X1 U1295 ( .A(n1334), .B(n1335), .C(n1336), .Y(n1329) );
  AND2X1 U1296 ( .A(n1337), .B(n1338), .Y(n1336) );
  OAI21X1 U1297 ( .A(n1339), .B(n1340), .C(n1341), .Y(n1335) );
  AOI21X1 U1298 ( .A(n1342), .B(n1343), .C(n1344), .Y(n1340) );
  OAI21X1 U1299 ( .A(n1345), .B(n1346), .C(n1347), .Y(n1342) );
  AOI21X1 U1300 ( .A(n1348), .B(n1349), .C(n1350), .Y(n1346) );
  NAND2X1 U1301 ( .A(n1351), .B(n1352), .Y(n1350) );
  OAI21X1 U1302 ( .A(n1353), .B(n1354), .C(n1355), .Y(n1348) );
  AOI21X1 U1303 ( .A(n1356), .B(n1357), .C(n1358), .Y(n1354) );
  OAI21X1 U1304 ( .A(n1359), .B(n1360), .C(n1361), .Y(n1356) );
  AOI21X1 U1305 ( .A(n1362), .B(n1363), .C(n1364), .Y(n1360) );
  OAI21X1 U1306 ( .A(n1365), .B(n1366), .C(n1367), .Y(n1363) );
  NAND2X1 U1307 ( .A(n1368), .B(n1369), .Y(n1366) );
  AOI21X1 U1308 ( .A(n1370), .B(n1371), .C(n1372), .Y(n1365) );
  OAI21X1 U1309 ( .A(n1373), .B(n1374), .C(n1375), .Y(n1371) );
  OAI21X1 U1310 ( .A(n1376), .B(n1377), .C(n1378), .Y(n1374) );
  NAND2X1 U1311 ( .A(n1379), .B(n1380), .Y(n1377) );
  AOI21X1 U1312 ( .A(n1381), .B(n1382), .C(n1383), .Y(n1376) );
  OAI21X1 U1313 ( .A(n1384), .B(n1385), .C(n1386), .Y(n1381) );
  AOI21X1 U1314 ( .A(n1387), .B(n1388), .C(n1389), .Y(n1384) );
  INVX1 U1315 ( .A(n1390), .Y(n1389) );
  OAI21X1 U1316 ( .A(n1391), .B(n1392), .C(n1393), .Y(n1388) );
  AND2X1 U1317 ( .A(n1394), .B(n1395), .Y(n1391) );
  OAI21X1 U1318 ( .A(n1396), .B(n1397), .C(n1398), .Y(n1395) );
  OAI21X1 U1319 ( .A(n1399), .B(n1400), .C(n1401), .Y(n1397) );
  OAI21X1 U1320 ( .A(n1402), .B(n1403), .C(n1404), .Y(n1400) );
  AOI21X1 U1321 ( .A(n1405), .B(n1406), .C(n1407), .Y(n1402) );
  OAI21X1 U1322 ( .A(n1408), .B(n1409), .C(n1410), .Y(n1405) );
  AOI21X1 U1323 ( .A(n1411), .B(n1412), .C(n1413), .Y(n1409) );
  NAND3X1 U1324 ( .A(n1414), .B(n1415), .C(n1416), .Y(n1412) );
  OAI21X1 U1325 ( .A(n1417), .B(n1418), .C(n1419), .Y(n1411) );
  INVX1 U1326 ( .A(n1420), .Y(n1418) );
  AOI21X1 U1327 ( .A(n1421), .B(n1422), .C(n1423), .Y(n1417) );
  OAI21X1 U1328 ( .A(n1424), .B(n1425), .C(n1426), .Y(n1422) );
  AOI21X1 U1329 ( .A(n1427), .B(n1428), .C(n1429), .Y(n1424) );
  OAI21X1 U1330 ( .A(n1430), .B(n1431), .C(n1432), .Y(n1428) );
  AND2X1 U1331 ( .A(n1433), .B(n1434), .Y(n1432) );
  AOI21X1 U1332 ( .A(n1435), .B(n1436), .C(n1437), .Y(n1430) );
  INVX1 U1333 ( .A(n1438), .Y(n1437) );
  OAI21X1 U1334 ( .A(n1439), .B(n1440), .C(n1441), .Y(n1435) );
  OAI21X1 U1335 ( .A(n1442), .B(n1443), .C(n1444), .Y(n1440) );
  AOI22X1 U1336 ( .A(n1445), .B(n1446), .C(n1447), .D(n1448), .Y(n1443) );
  OAI22X1 U1337 ( .A(n1449), .B(n1258), .C(n1450), .D(n1451), .Y(n1445) );
  AOI22X1 U1338 ( .A(n1452), .B(n1453), .C(n1454), .D(n1455), .Y(n1450) );
  AND2X1 U1339 ( .A(n1456), .B(n1457), .Y(n1452) );
  INVX1 U1340 ( .A(n1458), .Y(n1449) );
  NAND2X1 U1341 ( .A(n1459), .B(n1460), .Y(n1396) );
  AND2X1 U1342 ( .A(n1461), .B(n1462), .Y(n1387) );
  NAND2X1 U1343 ( .A(n1463), .B(n1464), .Y(n1373) );
  INVX1 U1344 ( .A(n1465), .Y(n1370) );
  AND2X1 U1345 ( .A(n1466), .B(n1467), .Y(n1362) );
  INVX1 U1346 ( .A(n1468), .Y(n1359) );
  INVX1 U1347 ( .A(n1469), .Y(n1345) );
  INVX1 U1348 ( .A(n1470), .Y(n1300) );
  NAND2X1 U1349 ( .A(n1471), .B(n1472), .Y(n1274) );
  NAND2X1 U1350 ( .A(n1473), .B(n1474), .Y(n1268) );
  MUX2X1 U1351 ( .B(n1475), .A(n1476), .S(n1259), .Y(n1246) );
  OAI21X1 U1352 ( .A(n1477), .B(n1478), .C(n1479), .Y(n1475) );
  AOI21X1 U1353 ( .A(n1480), .B(n1481), .C(n1482), .Y(n1477) );
  INVX1 U1354 ( .A(n1483), .Y(n1482) );
  OAI21X1 U1355 ( .A(n1484), .B(n1485), .C(n1270), .Y(n1481) );
  AOI21X1 U1356 ( .A(n1273), .B(n1486), .C(n1487), .Y(n1484) );
  INVX1 U1357 ( .A(n1488), .Y(n1487) );
  NAND3X1 U1358 ( .A(n1489), .B(n1471), .C(n1278), .Y(n1486) );
  OAI21X1 U1359 ( .A(n1490), .B(n1491), .C(n1281), .Y(n1489) );
  AOI21X1 U1360 ( .A(n1492), .B(n1493), .C(n1494), .Y(n1491) );
  INVX1 U1361 ( .A(n1495), .Y(n1494) );
  OAI21X1 U1362 ( .A(n1496), .B(n1497), .C(n1287), .Y(n1492) );
  AOI22X1 U1363 ( .A(n1498), .B(n1499), .C(n1500), .D(n1501), .Y(n1497) );
  OAI21X1 U1364 ( .A(n1502), .B(n1503), .C(n1504), .Y(n1499) );
  AOI21X1 U1365 ( .A(n1505), .B(n1506), .C(n1507), .Y(n1503) );
  OAI21X1 U1366 ( .A(n1508), .B(n1509), .C(n1299), .Y(n1506) );
  AOI21X1 U1367 ( .A(n1510), .B(n1511), .C(n1512), .Y(n1508) );
  NAND2X1 U1368 ( .A(n1513), .B(n1514), .Y(n1512) );
  OAI21X1 U1369 ( .A(n1515), .B(n1516), .C(n1517), .Y(n1511) );
  INVX1 U1370 ( .A(n1308), .Y(n1517) );
  AOI21X1 U1371 ( .A(n1518), .B(n1322), .C(n1519), .Y(n1516) );
  NAND3X1 U1372 ( .A(n1520), .B(n1521), .C(n1522), .Y(n1518) );
  AOI22X1 U1373 ( .A(n1523), .B(n1524), .C(n1525), .D(n1526), .Y(n1522) );
  AOI21X1 U1374 ( .A(n1325), .B(n1527), .C(n1528), .Y(n1523) );
  INVX1 U1375 ( .A(n1529), .Y(n1528) );
  OAI21X1 U1376 ( .A(n1530), .B(n1531), .C(n1532), .Y(n1527) );
  AND2X1 U1377 ( .A(n1533), .B(n1534), .Y(n1532) );
  AOI21X1 U1378 ( .A(n1535), .B(n1536), .C(n1537), .Y(n1530) );
  NAND2X1 U1379 ( .A(n1538), .B(n1338), .Y(n1537) );
  OAI21X1 U1380 ( .A(n1539), .B(n1540), .C(n1541), .Y(n1536) );
  AOI21X1 U1381 ( .A(n1542), .B(n1543), .C(n1344), .Y(n1540) );
  INVX1 U1382 ( .A(n1544), .Y(n1344) );
  OAI21X1 U1383 ( .A(n1545), .B(n1546), .C(n1547), .Y(n1542) );
  AOI21X1 U1384 ( .A(n1548), .B(n1357), .C(n1549), .Y(n1545) );
  NAND2X1 U1385 ( .A(n1550), .B(n1551), .Y(n1549) );
  OAI21X1 U1386 ( .A(n1552), .B(n1553), .C(n1554), .Y(n1548) );
  AND2X1 U1387 ( .A(n1555), .B(n1468), .Y(n1554) );
  AOI21X1 U1388 ( .A(n1556), .B(n1557), .C(n1364), .Y(n1552) );
  OAI21X1 U1389 ( .A(n1558), .B(n1559), .C(n1367), .Y(n1557) );
  INVX1 U1390 ( .A(n1368), .Y(n1559) );
  AOI21X1 U1391 ( .A(n1560), .B(n1561), .C(n1562), .Y(n1558) );
  AOI21X1 U1392 ( .A(n1563), .B(n1564), .C(n1465), .Y(n1560) );
  OAI21X1 U1393 ( .A(n1565), .B(n1566), .C(n1567), .Y(n1465) );
  OAI21X1 U1394 ( .A(n1568), .B(n1569), .C(n1570), .Y(n1564) );
  AOI21X1 U1395 ( .A(n1571), .B(n1378), .C(n1572), .Y(n1569) );
  INVX1 U1396 ( .A(n1379), .Y(n1572) );
  NAND3X1 U1397 ( .A(n1573), .B(n1574), .C(n1575), .Y(n1571) );
  OAI21X1 U1398 ( .A(n1576), .B(n1577), .C(n1578), .Y(n1575) );
  AND2X1 U1399 ( .A(n1579), .B(n1380), .Y(n1578) );
  AOI21X1 U1400 ( .A(n1580), .B(n1581), .C(n1582), .Y(n1577) );
  OAI21X1 U1401 ( .A(n1583), .B(n1584), .C(n1585), .Y(n1580) );
  OAI21X1 U1402 ( .A(n1586), .B(n1587), .C(n1588), .Y(n1584) );
  NAND2X1 U1403 ( .A(n1589), .B(n1393), .Y(n1587) );
  AOI21X1 U1404 ( .A(n1590), .B(n1591), .C(n1592), .Y(n1586) );
  OAI21X1 U1405 ( .A(n1593), .B(n1594), .C(n1595), .Y(n1590) );
  AOI21X1 U1406 ( .A(n1596), .B(n1401), .C(n1597), .Y(n1594) );
  OAI21X1 U1407 ( .A(n1598), .B(n1599), .C(n1600), .Y(n1596) );
  NAND3X1 U1408 ( .A(n1416), .B(n1601), .C(n1602), .Y(n1600) );
  AOI21X1 U1409 ( .A(n1603), .B(n1604), .C(n1605), .Y(n1598) );
  INVX1 U1410 ( .A(n1404), .Y(n1605) );
  OAI21X1 U1411 ( .A(n1606), .B(n1607), .C(n1608), .Y(n1604) );
  NAND2X1 U1412 ( .A(n1406), .B(n1609), .Y(n1607) );
  AOI21X1 U1413 ( .A(n1610), .B(n1611), .C(n1612), .Y(n1606) );
  OAI21X1 U1414 ( .A(n1613), .B(n1614), .C(n1615), .Y(n1610) );
  AOI21X1 U1415 ( .A(n1426), .B(n1616), .C(n1617), .Y(n1614) );
  OAI21X1 U1416 ( .A(n1429), .B(n1618), .C(n1619), .Y(n1616) );
  AOI21X1 U1417 ( .A(n1620), .B(n1621), .C(n1622), .Y(n1618) );
  OAI21X1 U1418 ( .A(n1623), .B(n1624), .C(n1625), .Y(n1620) );
  OAI21X1 U1419 ( .A(n1442), .B(n1626), .C(n1627), .Y(n1624) );
  OAI21X1 U1420 ( .A(n1628), .B(n1629), .C(n1630), .Y(n1627) );
  AOI21X1 U1421 ( .A(n1458), .B(n1476), .C(n1631), .Y(n1626) );
  NAND3X1 U1422 ( .A(n1632), .B(n1633), .C(n1455), .Y(n1458) );
  INVX1 U1423 ( .A(n1634), .Y(n1442) );
  NAND3X1 U1424 ( .A(n1447), .B(n1453), .C(n1635), .Y(n1634) );
  NOR2X1 U1425 ( .A(n1636), .B(n1637), .Y(n1635) );
  INVX1 U1426 ( .A(n1638), .Y(n1426) );
  NAND2X1 U1427 ( .A(n1639), .B(n1640), .Y(n1583) );
  NOR2X1 U1428 ( .A(n1641), .B(n1642), .Y(n1563) );
  INVX1 U1429 ( .A(n1643), .Y(n1515) );
  NOR2X1 U1430 ( .A(n1644), .B(n1645), .Y(n1498) );
  NAND2X1 U1431 ( .A(n1646), .B(n1647), .Y(n1244) );
  MUX2X1 U1432 ( .B(n1648), .A(state[3]), .S(n1259), .Y(n1646) );
  AOI22X1 U1433 ( .A(n1649), .B(n1650), .C(n1651), .D(n1652), .Y(n1648) );
  OAI21X1 U1434 ( .A(n1653), .B(n1260), .C(n1480), .Y(n1651) );
  AOI21X1 U1435 ( .A(n1654), .B(n1655), .C(n1267), .Y(n1653) );
  OAI21X1 U1436 ( .A(n1656), .B(n1657), .C(n1658), .Y(n1655) );
  OAI21X1 U1437 ( .A(n1659), .B(n1660), .C(n1661), .Y(n1657) );
  NAND2X1 U1438 ( .A(n1662), .B(n1663), .Y(n1661) );
  OAI21X1 U1439 ( .A(n1276), .B(n1664), .C(n1665), .Y(n1662) );
  OAI21X1 U1440 ( .A(n1666), .B(n1667), .C(n1668), .Y(n1664) );
  AOI21X1 U1441 ( .A(n1669), .B(n1670), .C(n1671), .Y(n1666) );
  NAND3X1 U1442 ( .A(n1504), .B(n1289), .C(n1672), .Y(n1670) );
  AOI21X1 U1443 ( .A(n1673), .B(n1674), .C(n1675), .Y(n1672) );
  AND2X1 U1444 ( .A(n1505), .B(n1676), .Y(n1674) );
  NAND3X1 U1445 ( .A(n1677), .B(n1678), .C(n1679), .Y(n1505) );
  AOI21X1 U1446 ( .A(n1680), .B(n1681), .C(n1682), .Y(n1673) );
  OAI21X1 U1447 ( .A(n1683), .B(n1684), .C(n1685), .Y(n1680) );
  AOI21X1 U1448 ( .A(n1686), .B(n1687), .C(n1509), .Y(n1684) );
  INVX1 U1449 ( .A(n1688), .Y(n1509) );
  NAND3X1 U1450 ( .A(n1513), .B(n1470), .C(n1689), .Y(n1686) );
  OAI21X1 U1451 ( .A(n1308), .B(n1690), .C(n1691), .Y(n1689) );
  NOR2X1 U1452 ( .A(n1692), .B(n1693), .Y(n1691) );
  OAI21X1 U1453 ( .A(n1694), .B(n1695), .C(n1313), .Y(n1690) );
  NAND2X1 U1454 ( .A(n1314), .B(n1696), .Y(n1695) );
  AOI21X1 U1455 ( .A(n1643), .B(n1697), .C(n1698), .Y(n1694) );
  NAND3X1 U1456 ( .A(n1520), .B(n1521), .C(n1699), .Y(n1697) );
  AOI21X1 U1457 ( .A(n1524), .B(n1700), .C(n1701), .Y(n1699) );
  OAI21X1 U1458 ( .A(n1531), .B(n1702), .C(n1703), .Y(n1700) );
  NAND3X1 U1459 ( .A(n1704), .B(n1705), .C(n1706), .Y(n1703) );
  AOI21X1 U1460 ( .A(n1707), .B(n1708), .C(n1709), .Y(n1702) );
  NAND2X1 U1461 ( .A(n1338), .B(n1710), .Y(n1709) );
  INVX1 U1462 ( .A(n1711), .Y(n1710) );
  OAI21X1 U1463 ( .A(n1712), .B(n1713), .C(n1714), .Y(n1708) );
  NAND2X1 U1464 ( .A(n1715), .B(n1343), .Y(n1713) );
  OAI21X1 U1465 ( .A(n1716), .B(n1717), .C(n1351), .Y(n1715) );
  INVX1 U1466 ( .A(n1718), .Y(n1717) );
  AOI21X1 U1467 ( .A(n1550), .B(n1719), .C(n1720), .Y(n1716) );
  OAI21X1 U1468 ( .A(n1721), .B(n1353), .C(n1349), .Y(n1719) );
  INVX1 U1469 ( .A(n1722), .Y(n1353) );
  AOI21X1 U1470 ( .A(n1723), .B(n1724), .C(n1725), .Y(n1721) );
  INVX1 U1471 ( .A(n1361), .Y(n1725) );
  OAI21X1 U1472 ( .A(n1726), .B(n1727), .C(n1728), .Y(n1724) );
  INVX1 U1473 ( .A(n1729), .Y(n1727) );
  AOI21X1 U1474 ( .A(n1730), .B(n1731), .C(n1732), .Y(n1726) );
  OAI21X1 U1475 ( .A(n1733), .B(n1734), .C(n1368), .Y(n1731) );
  AOI21X1 U1476 ( .A(n1735), .B(n1736), .C(n1737), .Y(n1733) );
  OAI21X1 U1477 ( .A(n1738), .B(n1739), .C(n1375), .Y(n1736) );
  NAND2X1 U1478 ( .A(n1740), .B(n1463), .Y(n1739) );
  AOI21X1 U1479 ( .A(n1379), .B(n1741), .C(n1568), .Y(n1738) );
  INVX1 U1480 ( .A(n1742), .Y(n1568) );
  NAND3X1 U1481 ( .A(n1573), .B(n1378), .C(n1743), .Y(n1741) );
  OAI21X1 U1482 ( .A(n1744), .B(n1745), .C(n1380), .Y(n1743) );
  AOI21X1 U1483 ( .A(n1382), .B(n1746), .C(n1747), .Y(n1744) );
  INVX1 U1484 ( .A(n1748), .Y(n1747) );
  OAI21X1 U1485 ( .A(n1749), .B(n1750), .C(n1581), .Y(n1746) );
  OAI22X1 U1486 ( .A(n1751), .B(n1752), .C(n1753), .D(n1754), .Y(n1750) );
  OAI21X1 U1487 ( .A(n1755), .B(n1756), .C(n1589), .Y(n1754) );
  AOI21X1 U1488 ( .A(n1757), .B(n1758), .C(n1759), .Y(n1756) );
  INVX1 U1489 ( .A(n1760), .Y(n1759) );
  AOI21X1 U1490 ( .A(n1761), .B(n1762), .C(n1763), .Y(n1757) );
  OAI21X1 U1491 ( .A(n1764), .B(n1765), .C(n1766), .Y(n1762) );
  AOI21X1 U1492 ( .A(n1767), .B(n1768), .C(n1769), .Y(n1764) );
  OAI21X1 U1493 ( .A(n1413), .B(n1770), .C(n1771), .Y(n1769) );
  OAI21X1 U1494 ( .A(n1772), .B(n1423), .C(n1611), .Y(n1770) );
  AOI21X1 U1495 ( .A(n1773), .B(n1774), .C(n1613), .Y(n1772) );
  INVX1 U1496 ( .A(n1775), .Y(n1613) );
  OAI21X1 U1497 ( .A(n1776), .B(n1777), .C(n1778), .Y(n1774) );
  AOI21X1 U1498 ( .A(n1779), .B(n1427), .C(n1429), .Y(n1777) );
  INVX1 U1499 ( .A(n1780), .Y(n1429) );
  OAI21X1 U1500 ( .A(n1622), .B(n1781), .C(n1434), .Y(n1779) );
  INVX1 U1501 ( .A(n1782), .Y(n1781) );
  OAI21X1 U1502 ( .A(n1783), .B(n1784), .C(n1621), .Y(n1782) );
  AOI21X1 U1503 ( .A(n1438), .B(n1785), .C(n1431), .Y(n1784) );
  OAI21X1 U1504 ( .A(n1786), .B(n1787), .C(n1788), .Y(n1431) );
  OR2X1 U1505 ( .A(n1789), .B(n1790), .Y(n1787) );
  NAND2X1 U1506 ( .A(n1791), .B(n1414), .Y(n1786) );
  INVX1 U1507 ( .A(n1792), .Y(n1785) );
  AOI21X1 U1508 ( .A(n1793), .B(n1794), .C(n1795), .Y(n1792) );
  OAI21X1 U1509 ( .A(n1796), .B(n1628), .C(n1630), .Y(n1794) );
  NOR2X1 U1510 ( .A(state[3]), .B(n1797), .Y(n1793) );
  INVX1 U1511 ( .A(n1798), .Y(n1622) );
  NOR2X1 U1512 ( .A(n1799), .B(n1800), .Y(n1767) );
  AND2X1 U1513 ( .A(n1801), .B(n1802), .Y(n1761) );
  OAI21X1 U1514 ( .A(n1803), .B(n1804), .C(n1805), .Y(n1801) );
  INVX1 U1515 ( .A(n1806), .Y(n1753) );
  NAND3X1 U1516 ( .A(n1639), .B(n1640), .C(n1585), .Y(n1749) );
  INVX1 U1517 ( .A(n1334), .Y(n1707) );
  NAND2X1 U1518 ( .A(n1488), .B(n1474), .Y(n1656) );
  NOR2X1 U1519 ( .A(n1799), .B(n1807), .Y(n1649) );
  NAND2X1 U1520 ( .A(n1808), .B(n1647), .Y(n1242) );
  MUX2X1 U1521 ( .B(n1809), .A(state[7]), .S(n1259), .Y(n1808) );
  AOI21X1 U1522 ( .A(n1479), .B(n1810), .C(n1811), .Y(n1809) );
  OAI21X1 U1523 ( .A(n1812), .B(n1264), .C(n1483), .Y(n1810) );
  NAND3X1 U1524 ( .A(n1813), .B(n1814), .C(n1704), .Y(n1483) );
  AOI21X1 U1525 ( .A(n1815), .B(n1816), .C(n1260), .Y(n1812) );
  OAI21X1 U1526 ( .A(n1817), .B(n1818), .C(n1270), .Y(n1816) );
  INVX1 U1527 ( .A(n1654), .Y(n1818) );
  AOI21X1 U1528 ( .A(n1273), .B(n1819), .C(n1485), .Y(n1817) );
  NAND2X1 U1529 ( .A(n1820), .B(n1473), .Y(n1819) );
  OAI21X1 U1530 ( .A(n1821), .B(n1822), .C(n1663), .Y(n1820) );
  AOI21X1 U1531 ( .A(n1823), .B(n1824), .C(n1825), .Y(n1822) );
  INVX1 U1532 ( .A(n1281), .Y(n1825) );
  OAI21X1 U1533 ( .A(n1667), .B(n1826), .C(n1827), .Y(n1823) );
  AOI21X1 U1534 ( .A(n1828), .B(n1293), .C(n1645), .Y(n1826) );
  INVX1 U1535 ( .A(n1288), .Y(n1645) );
  NAND3X1 U1536 ( .A(n1829), .B(n1633), .C(n1632), .Y(n1288) );
  OAI21X1 U1537 ( .A(n1830), .B(n1831), .C(n1832), .Y(n1828) );
  AOI21X1 U1538 ( .A(n1833), .B(n1685), .C(n1834), .Y(n1831) );
  NAND2X1 U1539 ( .A(n1681), .B(n1302), .Y(n1834) );
  OAI21X1 U1540 ( .A(n1835), .B(n1836), .C(n1837), .Y(n1833) );
  AOI21X1 U1541 ( .A(n1838), .B(n1314), .C(n1839), .Y(n1836) );
  OAI21X1 U1542 ( .A(n1840), .B(n1841), .C(n1842), .Y(n1838) );
  AOI21X1 U1543 ( .A(n1843), .B(n1322), .C(n1844), .Y(n1840) );
  OAI21X1 U1544 ( .A(n1845), .B(n1319), .C(n1846), .Y(n1843) );
  AND2X1 U1545 ( .A(n1323), .B(n1520), .Y(n1846) );
  NAND2X1 U1546 ( .A(n1521), .B(n1529), .Y(n1319) );
  NAND3X1 U1547 ( .A(n1847), .B(n1848), .C(n1849), .Y(n1529) );
  AOI21X1 U1548 ( .A(n1850), .B(n1328), .C(n1851), .Y(n1845) );
  OAI21X1 U1549 ( .A(n1852), .B(n1853), .C(n1854), .Y(n1850) );
  OAI21X1 U1550 ( .A(n1855), .B(n1856), .C(n1332), .Y(n1853) );
  OAI21X1 U1551 ( .A(n1857), .B(n1858), .C(n1338), .Y(n1856) );
  OAI21X1 U1552 ( .A(n1859), .B(n1860), .C(n1535), .Y(n1858) );
  NAND2X1 U1553 ( .A(n1544), .B(n1861), .Y(n1860) );
  AOI21X1 U1554 ( .A(n1862), .B(n1718), .C(n1863), .Y(n1859) );
  OAI21X1 U1555 ( .A(n1864), .B(n1865), .C(n1866), .Y(n1862) );
  AND2X1 U1556 ( .A(n1352), .B(n1543), .Y(n1866) );
  AOI21X1 U1557 ( .A(n1867), .B(n1868), .C(n1358), .Y(n1865) );
  OAI21X1 U1558 ( .A(n1869), .B(n1870), .C(n1871), .Y(n1868) );
  AND2X1 U1559 ( .A(n1872), .B(n1873), .Y(n1871) );
  AOI21X1 U1560 ( .A(n1729), .B(n1874), .C(n1364), .Y(n1869) );
  NAND3X1 U1561 ( .A(n1467), .B(n1466), .C(n1875), .Y(n1874) );
  OAI21X1 U1562 ( .A(n1876), .B(n1877), .C(n1556), .Y(n1875) );
  AOI21X1 U1563 ( .A(n1878), .B(n1368), .C(n1879), .Y(n1877) );
  OAI21X1 U1564 ( .A(n1880), .B(n1881), .C(n1882), .Y(n1878) );
  NOR2X1 U1565 ( .A(n1737), .B(n1734), .Y(n1882) );
  INVX1 U1566 ( .A(n1369), .Y(n1737) );
  AOI21X1 U1567 ( .A(n1883), .B(n1884), .C(n1885), .Y(n1880) );
  OAI21X1 U1568 ( .A(n1886), .B(n1887), .C(n1379), .Y(n1884) );
  OAI21X1 U1569 ( .A(n1888), .B(n1889), .C(n1378), .Y(n1887) );
  AOI21X1 U1570 ( .A(n1890), .B(n1891), .C(n1745), .Y(n1889) );
  INVX1 U1571 ( .A(n1892), .Y(n1745) );
  NAND3X1 U1572 ( .A(n1705), .B(n1633), .C(n1679), .Y(n1892) );
  OAI21X1 U1573 ( .A(n1893), .B(n1894), .C(n1581), .Y(n1891) );
  NAND3X1 U1574 ( .A(n1895), .B(n1678), .C(n1602), .Y(n1581) );
  AOI21X1 U1575 ( .A(n1896), .B(n1589), .C(n1897), .Y(n1894) );
  NAND2X1 U1576 ( .A(n1898), .B(n1461), .Y(n1897) );
  NAND2X1 U1577 ( .A(n1393), .B(n1899), .Y(n1896) );
  OAI21X1 U1578 ( .A(n1900), .B(n1901), .C(n1902), .Y(n1899) );
  NAND2X1 U1579 ( .A(n1394), .B(n1903), .Y(n1901) );
  OAI21X1 U1580 ( .A(n1904), .B(n1905), .C(n1906), .Y(n1903) );
  OAI21X1 U1581 ( .A(n1907), .B(n1908), .C(n1909), .Y(n1906) );
  OAI21X1 U1582 ( .A(n1910), .B(n1911), .C(n1398), .Y(n1908) );
  OAI21X1 U1583 ( .A(n1912), .B(n1913), .C(n1459), .Y(n1911) );
  NAND2X1 U1584 ( .A(n1802), .B(n1914), .Y(n1913) );
  NOR2X1 U1585 ( .A(n1407), .B(n1915), .Y(n1912) );
  INVX1 U1586 ( .A(n1916), .Y(n1915) );
  OAI21X1 U1587 ( .A(n1413), .B(n1917), .C(n1918), .Y(n1916) );
  OAI21X1 U1588 ( .A(n1919), .B(n1920), .C(n1406), .Y(n1917) );
  AOI21X1 U1589 ( .A(n1921), .B(n1775), .C(n1423), .Y(n1920) );
  NAND3X1 U1590 ( .A(n1922), .B(n1923), .C(n1924), .Y(n1775) );
  OAI21X1 U1591 ( .A(n1776), .B(n1925), .C(n1926), .Y(n1921) );
  AOI21X1 U1592 ( .A(n1927), .B(n1621), .C(n1928), .Y(n1925) );
  INVX1 U1593 ( .A(n1434), .Y(n1928) );
  NAND3X1 U1594 ( .A(n1796), .B(n1929), .C(n1930), .Y(n1621) );
  OAI21X1 U1595 ( .A(n1931), .B(n1623), .C(n1625), .Y(n1927) );
  AND2X1 U1596 ( .A(n1932), .B(n1438), .Y(n1625) );
  NAND2X1 U1597 ( .A(n1441), .B(n1788), .Y(n1623) );
  AOI21X1 U1598 ( .A(n1933), .B(n1444), .C(n1934), .Y(n1931) );
  INVX1 U1599 ( .A(n1935), .Y(n1934) );
  NOR2X1 U1600 ( .A(state[7]), .B(n1936), .Y(n1933) );
  INVX1 U1601 ( .A(n1419), .Y(n1919) );
  OAI21X1 U1602 ( .A(n1799), .B(n1937), .C(n1766), .Y(n1407) );
  NAND2X1 U1603 ( .A(n1938), .B(n1414), .Y(n1905) );
  INVX1 U1604 ( .A(n1632), .Y(n1904) );
  INVX1 U1605 ( .A(n1383), .Y(n1890) );
  NAND3X1 U1606 ( .A(n1579), .B(n1939), .C(n1748), .Y(n1383) );
  NAND3X1 U1607 ( .A(n1940), .B(n1414), .C(n1941), .Y(n1748) );
  NAND3X1 U1608 ( .A(n1416), .B(n1414), .C(n1940), .Y(n1579) );
  INVX1 U1609 ( .A(n1573), .Y(n1886) );
  NOR2X1 U1610 ( .A(n1641), .B(n1942), .Y(n1883) );
  INVX1 U1611 ( .A(n1367), .Y(n1876) );
  INVX1 U1612 ( .A(n1550), .Y(n1864) );
  INVX1 U1613 ( .A(n1943), .Y(n1857) );
  NAND2X1 U1614 ( .A(n1337), .B(n1330), .Y(n1855) );
  NAND2X1 U1615 ( .A(n1333), .B(n1533), .Y(n1852) );
  NAND3X1 U1616 ( .A(n1944), .B(n1601), .C(n1945), .Y(n1533) );
  INVX1 U1617 ( .A(n1687), .Y(n1835) );
  INVX1 U1618 ( .A(n1287), .Y(n1667) );
  INVX1 U1619 ( .A(n1946), .Y(n1821) );
  NAND2X1 U1620 ( .A(n1947), .B(n1948), .Y(n1240) );
  INVX1 U1621 ( .A(n1255), .Y(n1948) );
  OAI21X1 U1622 ( .A(n1949), .B(n1259), .C(n1647), .Y(n1255) );
  INVX1 U1623 ( .A(n1478), .Y(n1949) );
  AOI22X1 U1624 ( .A(n1950), .B(n1951), .C(state[6]), .D(n1259), .Y(n1947) );
  NOR2X1 U1625 ( .A(n1263), .B(n1260), .Y(n1951) );
  INVX1 U1626 ( .A(n1952), .Y(n1260) );
  AOI21X1 U1627 ( .A(n1953), .B(n1954), .C(n1955), .Y(n1950) );
  NAND3X1 U1628 ( .A(n1956), .B(n1488), .C(n1957), .Y(n1954) );
  OAI21X1 U1629 ( .A(n1958), .B(n1272), .C(n1273), .Y(n1957) );
  INVX1 U1630 ( .A(n1959), .Y(n1273) );
  AOI21X1 U1631 ( .A(n1960), .B(n1471), .C(n1961), .Y(n1958) );
  OAI21X1 U1632 ( .A(n1490), .B(n1962), .C(n1281), .Y(n1960) );
  NAND2X1 U1633 ( .A(n1963), .B(n1964), .Y(n1281) );
  AOI21X1 U1634 ( .A(n1965), .B(n1966), .C(n1967), .Y(n1962) );
  OAI21X1 U1635 ( .A(n1968), .B(n1969), .C(n1970), .Y(n1966) );
  NOR2X1 U1636 ( .A(n1644), .B(n1830), .Y(n1970) );
  INVX1 U1637 ( .A(n1289), .Y(n1644) );
  NAND2X1 U1638 ( .A(n1971), .B(n1676), .Y(n1969) );
  AOI21X1 U1639 ( .A(n1972), .B(n1973), .C(n1974), .Y(n1968) );
  NAND3X1 U1640 ( .A(n1513), .B(n1514), .C(n1975), .Y(n1973) );
  OAI21X1 U1641 ( .A(n1976), .B(n1977), .C(n1510), .Y(n1975) );
  NOR2X1 U1642 ( .A(n1978), .B(n1693), .Y(n1510) );
  AOI21X1 U1643 ( .A(n1979), .B(n1980), .C(n1981), .Y(n1977) );
  INVX1 U1644 ( .A(n1696), .Y(n1981) );
  NAND3X1 U1645 ( .A(n1982), .B(n1251), .C(n1938), .Y(n1696) );
  OAI21X1 U1646 ( .A(n1318), .B(n1983), .C(n1315), .Y(n1979) );
  AOI21X1 U1647 ( .A(n1984), .B(n1985), .C(n1844), .Y(n1983) );
  INVX1 U1648 ( .A(n1317), .Y(n1844) );
  NAND3X1 U1649 ( .A(n1986), .B(n1987), .C(n1988), .Y(n1317) );
  OAI21X1 U1650 ( .A(n1989), .B(n1990), .C(n1520), .Y(n1985) );
  AOI21X1 U1651 ( .A(n1991), .B(n1534), .C(n1851), .Y(n1989) );
  INVX1 U1652 ( .A(n1325), .Y(n1851) );
  OAI21X1 U1653 ( .A(n1326), .B(n1992), .C(n1854), .Y(n1991) );
  NAND3X1 U1654 ( .A(n1993), .B(n1982), .C(n1994), .Y(n1854) );
  AOI21X1 U1655 ( .A(n1995), .B(n1330), .C(n1996), .Y(n1992) );
  OAI21X1 U1656 ( .A(n1997), .B(n1334), .C(n1333), .Y(n1995) );
  NAND2X1 U1657 ( .A(n1538), .B(n1535), .Y(n1334) );
  AOI21X1 U1658 ( .A(n1998), .B(n1999), .C(n2000), .Y(n1997) );
  OAI21X1 U1659 ( .A(n1712), .B(n2001), .C(n1347), .Y(n1999) );
  OAI21X1 U1660 ( .A(n2002), .B(n2003), .C(n2004), .Y(n2001) );
  NOR2X1 U1661 ( .A(n1546), .B(n2005), .Y(n2003) );
  OAI21X1 U1662 ( .A(n2006), .B(n2007), .C(n2008), .Y(n2005) );
  OAI21X1 U1663 ( .A(n2009), .B(n2010), .C(n2011), .Y(n2008) );
  AND2X1 U1664 ( .A(n1550), .B(n1873), .Y(n2011) );
  OAI21X1 U1665 ( .A(n1553), .B(n2012), .C(n1468), .Y(n2010) );
  OAI21X1 U1666 ( .A(n2013), .B(n1732), .C(n1729), .Y(n2012) );
  NAND3X1 U1667 ( .A(n1804), .B(n1678), .C(n1988), .Y(n1729) );
  AOI21X1 U1668 ( .A(n2014), .B(n2015), .C(n2016), .Y(n2013) );
  NAND3X1 U1669 ( .A(n1561), .B(n2017), .C(n1735), .Y(n2015) );
  INVX1 U1670 ( .A(n2018), .Y(n1735) );
  NAND3X1 U1671 ( .A(n1567), .B(n2019), .C(n2020), .Y(n2018) );
  NAND2X1 U1672 ( .A(n2021), .B(n2022), .Y(n1567) );
  NAND3X1 U1673 ( .A(n1375), .B(n1464), .C(n2023), .Y(n2017) );
  OAI21X1 U1674 ( .A(n2024), .B(n2025), .C(n1378), .Y(n2023) );
  OAI21X1 U1675 ( .A(n2026), .B(n2027), .C(n2028), .Y(n2025) );
  NAND2X1 U1676 ( .A(n1386), .B(n1462), .Y(n2027) );
  NAND2X1 U1677 ( .A(n2029), .B(n2030), .Y(n1462) );
  AOI21X1 U1678 ( .A(n2031), .B(n1639), .C(n2032), .Y(n2026) );
  INVX1 U1679 ( .A(n1589), .Y(n2032) );
  OAI21X1 U1680 ( .A(n2033), .B(n1900), .C(n2034), .Y(n2031) );
  INVX1 U1681 ( .A(n2035), .Y(n1900) );
  AND2X1 U1682 ( .A(n1394), .B(n2036), .Y(n2033) );
  OAI21X1 U1683 ( .A(n1599), .B(n2037), .C(n1909), .Y(n2036) );
  OAI21X1 U1684 ( .A(n2038), .B(n2039), .C(n1459), .Y(n2037) );
  NAND2X1 U1685 ( .A(n1603), .B(n2040), .Y(n2039) );
  OAI21X1 U1686 ( .A(n2041), .B(n2042), .C(n1608), .Y(n2040) );
  AOI21X1 U1687 ( .A(n1963), .B(n2043), .C(n2044), .Y(n1608) );
  OAI21X1 U1688 ( .A(n2045), .B(n2046), .C(n2047), .Y(n2042) );
  INVX1 U1689 ( .A(n2048), .Y(n2047) );
  AOI21X1 U1690 ( .A(n2049), .B(n1615), .C(n1408), .Y(n2046) );
  OAI21X1 U1691 ( .A(n1423), .B(n2050), .C(n1419), .Y(n2049) );
  AOI21X1 U1692 ( .A(n2051), .B(n2052), .C(n2053), .Y(n2050) );
  OAI21X1 U1693 ( .A(n2054), .B(n2055), .C(n1773), .Y(n2051) );
  INVX1 U1694 ( .A(n1427), .Y(n2055) );
  NAND3X1 U1695 ( .A(n2056), .B(n2057), .C(n1526), .Y(n1427) );
  AOI21X1 U1696 ( .A(n1788), .B(n2058), .C(n1783), .Y(n2054) );
  OAI21X1 U1697 ( .A(n1439), .B(n2059), .C(n1441), .Y(n2058) );
  NAND2X1 U1698 ( .A(n2060), .B(n2061), .Y(n2059) );
  NAND3X1 U1699 ( .A(n1250), .B(n1414), .C(n1988), .Y(n1788) );
  NAND2X1 U1700 ( .A(n1609), .B(n2063), .Y(n2041) );
  INVX1 U1701 ( .A(n2064), .Y(n2063) );
  NAND2X1 U1702 ( .A(n1802), .B(n1404), .Y(n2038) );
  NAND2X1 U1703 ( .A(n2065), .B(n1460), .Y(n1599) );
  NAND3X1 U1704 ( .A(n2066), .B(n1677), .C(n2056), .Y(n1460) );
  NAND2X1 U1705 ( .A(n1585), .B(n1573), .Y(n2024) );
  AND2X1 U1706 ( .A(n2067), .B(n2068), .Y(n1561) );
  NOR2X1 U1707 ( .A(n1562), .B(n1879), .Y(n2014) );
  NAND2X1 U1708 ( .A(n2069), .B(n2070), .Y(n2007) );
  INVX1 U1709 ( .A(n1547), .Y(n2002) );
  INVX1 U1710 ( .A(n1701), .Y(n1984) );
  INVX1 U1711 ( .A(n2071), .Y(n1318) );
  INVX1 U1712 ( .A(n1314), .Y(n1976) );
  NAND3X1 U1713 ( .A(n1796), .B(n2072), .C(n2073), .Y(n1513) );
  NOR2X1 U1714 ( .A(n2074), .B(n2075), .Y(n1972) );
  AND2X1 U1715 ( .A(n1493), .B(n1287), .Y(n1965) );
  NOR2X1 U1716 ( .A(n2076), .B(n1485), .Y(n1953) );
  INVX1 U1717 ( .A(n1658), .Y(n1485) );
  MUX2X1 U1718 ( .B(n2077), .A(n2078), .S(n1259), .Y(n1238) );
  NAND2X1 U1719 ( .A(n2079), .B(n2080), .Y(n2077) );
  OAI21X1 U1720 ( .A(n2081), .B(n1263), .C(n1652), .Y(n2080) );
  AOI21X1 U1721 ( .A(n1658), .B(n2082), .C(n2083), .Y(n2081) );
  NAND2X1 U1722 ( .A(n1956), .B(n1480), .Y(n2083) );
  OAI21X1 U1723 ( .A(n2084), .B(n1959), .C(n1488), .Y(n2082) );
  NAND3X1 U1724 ( .A(n1986), .B(n2085), .C(n1679), .Y(n1488) );
  OAI21X1 U1725 ( .A(n1659), .B(n1660), .C(n2086), .Y(n1959) );
  INVX1 U1726 ( .A(n1448), .Y(n1660) );
  AOI21X1 U1727 ( .A(n1278), .B(n2087), .C(n2088), .Y(n2084) );
  INVX1 U1728 ( .A(n1473), .Y(n2088) );
  NAND2X1 U1729 ( .A(n1813), .B(n2089), .Y(n1473) );
  OAI21X1 U1730 ( .A(n1967), .B(n2090), .C(n2091), .Y(n2087) );
  AND2X1 U1731 ( .A(n1471), .B(n1824), .Y(n2091) );
  OAI21X1 U1732 ( .A(n2092), .B(n2093), .C(n1495), .Y(n2090) );
  NAND2X1 U1733 ( .A(n1287), .B(n1493), .Y(n2093) );
  AOI21X1 U1734 ( .A(n2094), .B(n2095), .C(n1496), .Y(n2092) );
  NAND3X1 U1735 ( .A(n1676), .B(n1289), .C(n2096), .Y(n2095) );
  OAI21X1 U1736 ( .A(n2097), .B(n1974), .C(n2098), .Y(n2096) );
  NOR2X1 U1737 ( .A(n1507), .B(n2074), .Y(n2098) );
  INVX1 U1738 ( .A(n1681), .Y(n2074) );
  AOI21X1 U1739 ( .A(n2099), .B(n1687), .C(n2100), .Y(n2097) );
  OAI21X1 U1740 ( .A(n1303), .B(n2101), .C(n1470), .Y(n2099) );
  NAND3X1 U1741 ( .A(n2085), .B(n1414), .C(n1945), .Y(n1470) );
  AOI21X1 U1742 ( .A(n2102), .B(n1310), .C(n1693), .Y(n2101) );
  INVX1 U1743 ( .A(n1692), .Y(n1310) );
  NOR2X1 U1744 ( .A(n2103), .B(n2104), .Y(n1692) );
  OAI21X1 U1745 ( .A(n1308), .B(n2105), .C(n1314), .Y(n2102) );
  NAND3X1 U1746 ( .A(n2066), .B(n1796), .C(n2106), .Y(n1314) );
  OAI21X1 U1747 ( .A(n2107), .B(n1841), .C(n1643), .Y(n2105) );
  NAND2X1 U1748 ( .A(n1980), .B(n2071), .Y(n1841) );
  AOI21X1 U1749 ( .A(n2108), .B(n2109), .C(n1701), .Y(n2107) );
  OAI21X1 U1750 ( .A(n2110), .B(n2111), .C(n1322), .Y(n1701) );
  NAND3X1 U1751 ( .A(n1848), .B(n2112), .C(n2113), .Y(n1322) );
  OAI21X1 U1752 ( .A(n2114), .B(n1996), .C(n1524), .Y(n2109) );
  INVX1 U1753 ( .A(n1990), .Y(n1524) );
  NAND2X1 U1754 ( .A(n1323), .B(n2115), .Y(n1990) );
  NAND3X1 U1755 ( .A(n2072), .B(n2116), .C(n2117), .Y(n1323) );
  NOR2X1 U1756 ( .A(n2104), .B(n2006), .Y(n2117) );
  INVX1 U1757 ( .A(n2118), .Y(n2006) );
  AOI21X1 U1758 ( .A(n1333), .B(n2119), .C(n1711), .Y(n2114) );
  NOR2X1 U1759 ( .A(n2103), .B(n2120), .Y(n1711) );
  NAND3X1 U1760 ( .A(n1629), .B(state[2]), .C(n2069), .Y(n2103) );
  NAND3X1 U1761 ( .A(n1538), .B(n1338), .C(n2121), .Y(n2119) );
  OAI21X1 U1762 ( .A(n2122), .B(n2123), .C(n1535), .Y(n2121) );
  AOI21X1 U1763 ( .A(n2124), .B(n1541), .C(n2125), .Y(n2123) );
  OAI21X1 U1764 ( .A(n1339), .B(n2126), .C(n1341), .Y(n2124) );
  NAND3X1 U1765 ( .A(n2127), .B(n1986), .C(n1940), .Y(n1341) );
  AOI21X1 U1766 ( .A(n2128), .B(n1343), .C(n2129), .Y(n2126) );
  OAI21X1 U1767 ( .A(n2130), .B(n1712), .C(n1347), .Y(n2128) );
  AOI21X1 U1768 ( .A(n1351), .B(n2131), .C(n1863), .Y(n2130) );
  INVX1 U1769 ( .A(n2004), .Y(n1863) );
  NAND3X1 U1770 ( .A(n1718), .B(n1352), .C(n2132), .Y(n2131) );
  OAI21X1 U1771 ( .A(n1358), .B(n2133), .C(n1722), .Y(n2132) );
  AOI21X1 U1772 ( .A(n2134), .B(n2135), .C(n2136), .Y(n2133) );
  NAND2X1 U1773 ( .A(n2137), .B(n1361), .Y(n2136) );
  OAI21X1 U1774 ( .A(n1364), .B(n2138), .C(n1728), .Y(n2135) );
  AOI21X1 U1775 ( .A(n2139), .B(n1556), .C(n1732), .Y(n2138) );
  INVX1 U1776 ( .A(n1466), .Y(n1732) );
  OAI21X1 U1777 ( .A(n1734), .B(n2140), .C(n1730), .Y(n2139) );
  AOI21X1 U1778 ( .A(n2141), .B(n2142), .C(n1562), .Y(n2140) );
  INVX1 U1779 ( .A(n2143), .Y(n1562) );
  NAND3X1 U1780 ( .A(n1848), .B(n1677), .C(n1930), .Y(n2143) );
  INVX1 U1781 ( .A(n1881), .Y(n2142) );
  AOI21X1 U1782 ( .A(n2020), .B(n2144), .C(n1372), .Y(n2141) );
  INVX1 U1783 ( .A(n2145), .Y(n1372) );
  OAI21X1 U1784 ( .A(n2146), .B(n1642), .C(n2147), .Y(n2144) );
  OAI21X1 U1785 ( .A(n2022), .B(n1796), .C(n2021), .Y(n2147) );
  INVX1 U1786 ( .A(n1375), .Y(n1642) );
  AND2X1 U1787 ( .A(n2148), .B(n1740), .Y(n2146) );
  OAI21X1 U1788 ( .A(n2149), .B(n2150), .C(n2067), .Y(n2148) );
  OAI21X1 U1789 ( .A(n2151), .B(n2152), .C(n2153), .Y(n2150) );
  OAI21X1 U1790 ( .A(n1888), .B(n2154), .C(n1573), .Y(n2152) );
  NAND2X1 U1791 ( .A(n2155), .B(n2156), .Y(n1573) );
  AOI21X1 U1792 ( .A(n2157), .B(n1386), .C(n1576), .Y(n2154) );
  INVX1 U1793 ( .A(n1382), .Y(n1576) );
  NAND2X1 U1794 ( .A(n2158), .B(n1963), .Y(n1382) );
  OAI21X1 U1795 ( .A(n2159), .B(n2160), .C(n2161), .Y(n2157) );
  OAI21X1 U1796 ( .A(n2162), .B(n2163), .C(n1588), .Y(n2161) );
  INVX1 U1797 ( .A(n2164), .Y(n2163) );
  OAI21X1 U1798 ( .A(n2165), .B(n2166), .C(n1393), .Y(n2164) );
  NAND3X1 U1799 ( .A(n1758), .B(n2167), .C(n2035), .Y(n2166) );
  NAND3X1 U1800 ( .A(n1603), .B(n2168), .C(n2169), .Y(n2167) );
  NOR2X1 U1801 ( .A(n1910), .B(n1593), .Y(n2169) );
  INVX1 U1802 ( .A(n2170), .Y(n1593) );
  INVX1 U1803 ( .A(n1401), .Y(n1910) );
  OAI21X1 U1804 ( .A(n2171), .B(n2172), .C(n2173), .Y(n2168) );
  OAI21X1 U1805 ( .A(n2174), .B(n2044), .C(n2175), .Y(n2173) );
  INVX1 U1806 ( .A(n1403), .Y(n2175) );
  NAND2X1 U1807 ( .A(n2176), .B(n1609), .Y(n1403) );
  NAND3X1 U1808 ( .A(n1988), .B(n1982), .C(n2030), .Y(n1609) );
  INVX1 U1809 ( .A(n1766), .Y(n2044) );
  NAND3X1 U1810 ( .A(n2177), .B(n2178), .C(n2179), .Y(n1766) );
  NOR2X1 U1811 ( .A(n1637), .B(n2159), .Y(n2179) );
  NOR2X1 U1812 ( .A(n2180), .B(n1636), .Y(n2177) );
  AOI21X1 U1813 ( .A(n2181), .B(n2182), .C(n2064), .Y(n2174) );
  NAND3X1 U1814 ( .A(n2183), .B(n1611), .C(n2184), .Y(n2182) );
  INVX1 U1815 ( .A(n1413), .Y(n2184) );
  OAI21X1 U1816 ( .A(n2185), .B(n2186), .C(n2187), .Y(n1413) );
  NAND2X1 U1817 ( .A(n1414), .B(n1415), .Y(n2186) );
  INVX1 U1818 ( .A(n1796), .Y(n2185) );
  OAI21X1 U1819 ( .A(n1423), .B(n2188), .C(n1420), .Y(n2183) );
  AOI21X1 U1820 ( .A(n2189), .B(n1773), .C(n2053), .Y(n2188) );
  OAI21X1 U1821 ( .A(n1425), .B(n2190), .C(n2191), .Y(n2189) );
  AOI21X1 U1822 ( .A(n2192), .B(n1434), .C(n1776), .Y(n2190) );
  INVX1 U1823 ( .A(n1619), .Y(n1776) );
  NAND3X1 U1824 ( .A(n1250), .B(n1501), .C(n1982), .Y(n1619) );
  NAND3X1 U1825 ( .A(n1944), .B(n2066), .C(n1930), .Y(n1434) );
  OAI21X1 U1826 ( .A(n2193), .B(n1783), .C(n1798), .Y(n2192) );
  NAND3X1 U1827 ( .A(n1416), .B(state[2]), .C(n2194), .Y(n1798) );
  NOR2X1 U1828 ( .A(n2195), .B(n2159), .Y(n2194) );
  AOI22X1 U1829 ( .A(n2196), .B(n2197), .C(n2198), .D(n1438), .Y(n2193) );
  NAND2X1 U1830 ( .A(n1963), .B(n2089), .Y(n1438) );
  OAI21X1 U1831 ( .A(n2199), .B(n2200), .C(n2201), .Y(n2198) );
  NOR2X1 U1832 ( .A(n1936), .B(n2202), .Y(n2201) );
  INVX1 U1833 ( .A(n2203), .Y(n1936) );
  NAND2X1 U1834 ( .A(n1935), .B(n2060), .Y(n2200) );
  NAND3X1 U1835 ( .A(n2204), .B(n1803), .C(n1986), .Y(n1935) );
  NAND2X1 U1836 ( .A(n1444), .B(n2078), .Y(n2199) );
  INVX1 U1837 ( .A(state[5]), .Y(n2078) );
  NAND2X1 U1838 ( .A(n1630), .B(n1251), .Y(n1444) );
  NOR2X1 U1839 ( .A(n1789), .B(n2205), .Y(n2196) );
  INVX1 U1840 ( .A(n1778), .Y(n1425) );
  INVX1 U1841 ( .A(n2206), .Y(n1423) );
  NOR2X1 U1842 ( .A(n1612), .B(n2207), .Y(n2181) );
  INVX1 U1843 ( .A(n1399), .Y(n1603) );
  OAI21X1 U1844 ( .A(n2208), .B(n2172), .C(n1914), .Y(n1399) );
  INVX1 U1845 ( .A(n1805), .Y(n2172) );
  NAND3X1 U1846 ( .A(n1398), .B(n2209), .C(n1595), .Y(n2165) );
  NAND2X1 U1847 ( .A(n1963), .B(n1814), .Y(n2160) );
  INVX1 U1848 ( .A(n1380), .Y(n1888) );
  NAND2X1 U1849 ( .A(n1940), .B(n1963), .Y(n1380) );
  NAND2X1 U1850 ( .A(n1574), .B(n1379), .Y(n2151) );
  NAND3X1 U1851 ( .A(n2210), .B(n1929), .C(n2030), .Y(n1379) );
  NAND3X1 U1852 ( .A(n1463), .B(n1464), .C(n1378), .Y(n2149) );
  INVX1 U1853 ( .A(n2211), .Y(n1734) );
  INVX1 U1854 ( .A(n2212), .Y(n1364) );
  INVX1 U1855 ( .A(n1553), .Y(n2134) );
  NAND2X1 U1856 ( .A(n1723), .B(n1872), .Y(n1553) );
  NAND3X1 U1857 ( .A(n2213), .B(n1803), .C(n1982), .Y(n1872) );
  INVX1 U1858 ( .A(n1551), .Y(n1358) );
  NAND3X1 U1859 ( .A(n1796), .B(n2213), .C(n1633), .Y(n1352) );
  NAND3X1 U1860 ( .A(n2085), .B(n2214), .C(n1922), .Y(n1718) );
  NAND3X1 U1861 ( .A(n1922), .B(n1704), .C(n1849), .Y(n1351) );
  INVX1 U1862 ( .A(n2215), .Y(n2122) );
  NAND3X1 U1863 ( .A(n1601), .B(n1677), .C(n1993), .Y(n1338) );
  AND2X1 U1864 ( .A(n1521), .B(n1520), .Y(n2108) );
  INVX1 U1865 ( .A(n1514), .Y(n1303) );
  NOR2X1 U1866 ( .A(n2216), .B(n1671), .Y(n2094) );
  INVX1 U1867 ( .A(n2217), .Y(n1671) );
  NAND3X1 U1868 ( .A(n1964), .B(n1982), .C(n2218), .Y(n2217) );
  OAI21X1 U1869 ( .A(n2219), .B(n2220), .C(n1668), .Y(n1967) );
  NAND2X1 U1870 ( .A(n1628), .B(n1704), .Y(n2220) );
  NAND2X1 U1871 ( .A(n1414), .B(n2221), .Y(n2219) );
  INVX1 U1872 ( .A(n1961), .Y(n1278) );
  OAI21X1 U1873 ( .A(n2222), .B(n1955), .C(n2223), .Y(n1236) );
  INVX1 U1874 ( .A(n2224), .Y(n2223) );
  MUX2X1 U1875 ( .B(n2079), .A(n2225), .S(n1259), .Y(n2224) );
  NOR2X1 U1876 ( .A(n1811), .B(n1267), .Y(n2079) );
  INVX1 U1877 ( .A(n1815), .Y(n1267) );
  INVX1 U1878 ( .A(n2226), .Y(n1811) );
  NAND3X1 U1879 ( .A(n2227), .B(n1476), .C(n2113), .Y(n2226) );
  AOI21X1 U1880 ( .A(n2228), .B(n2229), .C(n1478), .Y(n2222) );
  NOR2X1 U1881 ( .A(n1285), .B(n2230), .Y(n1478) );
  INVX1 U1882 ( .A(n1501), .Y(n1285) );
  OAI21X1 U1883 ( .A(n2231), .B(n2232), .C(n1654), .Y(n2229) );
  AOI21X1 U1884 ( .A(n1448), .B(n2089), .C(n2233), .Y(n2232) );
  OAI21X1 U1885 ( .A(n1272), .B(n2234), .C(n1658), .Y(n2233) );
  NAND3X1 U1886 ( .A(n2235), .B(n1848), .C(n2236), .Y(n1658) );
  AND2X1 U1887 ( .A(n1633), .B(n2085), .Y(n2236) );
  INVX1 U1888 ( .A(n2237), .Y(n1848) );
  AOI22X1 U1889 ( .A(n2238), .B(n1986), .C(n2239), .D(n1946), .Y(n2234) );
  NAND3X1 U1890 ( .A(n1471), .B(n2240), .C(n2241), .Y(n2239) );
  AOI21X1 U1891 ( .A(n2242), .B(n2243), .C(n2244), .Y(n2241) );
  OAI21X1 U1892 ( .A(n2245), .B(n2246), .C(n1827), .Y(n2243) );
  INVX1 U1893 ( .A(n1280), .Y(n1827) );
  NAND2X1 U1894 ( .A(n2247), .B(n1668), .Y(n1280) );
  NAND2X1 U1895 ( .A(n1293), .B(n1287), .Y(n2246) );
  NAND2X1 U1896 ( .A(n2248), .B(n2213), .Y(n1287) );
  AOI21X1 U1897 ( .A(n2249), .B(n1504), .C(n1292), .Y(n2245) );
  INVX1 U1898 ( .A(n1676), .Y(n1292) );
  NAND3X1 U1899 ( .A(n2250), .B(n1629), .C(n1986), .Y(n1676) );
  OAI21X1 U1900 ( .A(n1682), .B(n2251), .C(n2252), .Y(n2249) );
  NOR2X1 U1901 ( .A(n1502), .B(n1507), .Y(n2252) );
  INVX1 U1902 ( .A(n1971), .Y(n1507) );
  INVX1 U1903 ( .A(n1298), .Y(n1502) );
  AOI21X1 U1904 ( .A(n2253), .B(n2254), .C(n1295), .Y(n2251) );
  NAND2X1 U1905 ( .A(n1688), .B(n1685), .Y(n1295) );
  NAND3X1 U1906 ( .A(n1895), .B(n1704), .C(n2255), .Y(n1688) );
  NOR2X1 U1907 ( .A(n1637), .B(n2256), .Y(n2255) );
  OAI21X1 U1908 ( .A(n2075), .B(n2257), .C(n1687), .Y(n2254) );
  NAND3X1 U1909 ( .A(n2227), .B(state[1]), .C(n1963), .Y(n1687) );
  AOI21X1 U1910 ( .A(n2258), .B(n1306), .C(n1693), .Y(n2257) );
  INVX1 U1911 ( .A(n2259), .Y(n1693) );
  NAND3X1 U1912 ( .A(n1986), .B(n2022), .C(n2260), .Y(n2259) );
  OAI21X1 U1913 ( .A(n1978), .B(n2261), .C(n2262), .Y(n2258) );
  NAND3X1 U1914 ( .A(n1633), .B(n1796), .C(n1938), .Y(n2262) );
  AOI21X1 U1915 ( .A(n2263), .B(n1980), .C(n1308), .Y(n2261) );
  OAI21X1 U1916 ( .A(n2230), .B(n2264), .C(n2265), .Y(n1308) );
  NAND3X1 U1917 ( .A(n1982), .B(n1629), .C(n1938), .Y(n2265) );
  OAI21X1 U1918 ( .A(n2266), .B(n2267), .C(n2071), .Y(n2263) );
  NAND2X1 U1919 ( .A(n2260), .B(n2113), .Y(n2071) );
  OAI21X1 U1920 ( .A(n2268), .B(n2269), .C(n1520), .Y(n2267) );
  NAND2X1 U1921 ( .A(n1525), .B(n1632), .Y(n1520) );
  INVX1 U1922 ( .A(n2111), .Y(n1525) );
  AOI21X1 U1923 ( .A(n2270), .B(n1325), .C(n2271), .Y(n2269) );
  INVX1 U1924 ( .A(n1521), .Y(n2271) );
  NAND3X1 U1925 ( .A(n2089), .B(n1678), .C(n2272), .Y(n1521) );
  OAI21X1 U1926 ( .A(n2273), .B(n2274), .C(n1534), .Y(n2270) );
  NAND3X1 U1927 ( .A(n1941), .B(n2057), .C(n1930), .Y(n1534) );
  AOI21X1 U1928 ( .A(n2275), .B(n2276), .C(n1996), .Y(n2274) );
  INVX1 U1929 ( .A(n1332), .Y(n1996) );
  NAND3X1 U1930 ( .A(n1601), .B(n1791), .C(n2277), .Y(n1332) );
  NOR2X1 U1931 ( .A(n1790), .B(n2278), .Y(n2277) );
  INVX1 U1932 ( .A(n1636), .Y(n1791) );
  OAI21X1 U1933 ( .A(n2000), .B(n2279), .C(n1337), .Y(n2276) );
  AOI21X1 U1934 ( .A(n2280), .B(n1544), .C(n1339), .Y(n2279) );
  OAI21X1 U1935 ( .A(n2281), .B(n2282), .C(n1343), .Y(n2280) );
  AOI21X1 U1936 ( .A(n1543), .B(n2283), .C(n1712), .Y(n2281) );
  OAI21X1 U1937 ( .A(n2284), .B(n2285), .C(n1469), .Y(n1712) );
  NAND3X1 U1938 ( .A(n1829), .B(n1601), .C(n1895), .Y(n1469) );
  NAND2X1 U1939 ( .A(n2066), .B(n1804), .Y(n2285) );
  INVX1 U1940 ( .A(n1706), .Y(n2284) );
  OAI21X1 U1941 ( .A(n1546), .B(n2286), .C(n1547), .Y(n2283) );
  NAND3X1 U1942 ( .A(n2287), .B(n1678), .C(n2260), .Y(n1547) );
  OAI21X1 U1943 ( .A(n2288), .B(n2289), .C(n1722), .Y(n2286) );
  NAND2X1 U1944 ( .A(n2043), .B(n1813), .Y(n1722) );
  NAND2X1 U1945 ( .A(n1873), .B(n1550), .Y(n2289) );
  NAND2X1 U1946 ( .A(n2290), .B(n1940), .Y(n1550) );
  AOI21X1 U1947 ( .A(n2291), .B(n1361), .C(n2292), .Y(n2288) );
  NAND3X1 U1948 ( .A(n1501), .B(n1678), .C(n2022), .Y(n1361) );
  OAI21X1 U1949 ( .A(n1870), .B(n2293), .C(n1468), .Y(n2291) );
  AOI21X1 U1950 ( .A(n2294), .B(n2295), .C(n2009), .Y(n2293) );
  NAND2X1 U1951 ( .A(n1728), .B(n1555), .Y(n2009) );
  NAND3X1 U1952 ( .A(n2250), .B(n1414), .C(n1803), .Y(n1555) );
  OAI21X1 U1953 ( .A(n1879), .B(n2296), .C(n1367), .Y(n2295) );
  NAND3X1 U1954 ( .A(n1945), .B(n1944), .C(n1986), .Y(n1367) );
  NOR2X1 U1955 ( .A(n2297), .B(n2298), .Y(n2296) );
  OAI21X1 U1956 ( .A(n1881), .B(n2299), .C(n2020), .Y(n2298) );
  OAI21X1 U1957 ( .A(n2300), .B(n2301), .C(n1375), .Y(n2299) );
  NAND3X1 U1958 ( .A(n1704), .B(n1250), .C(n1930), .Y(n1375) );
  INVX1 U1959 ( .A(n1740), .Y(n2301) );
  AOI21X1 U1960 ( .A(n2302), .B(n2303), .C(n1885), .Y(n2300) );
  INVX1 U1961 ( .A(n2067), .Y(n1885) );
  NAND2X1 U1962 ( .A(n2043), .B(n2248), .Y(n2067) );
  AND2X1 U1963 ( .A(n1464), .B(n1463), .Y(n2303) );
  NAND2X1 U1964 ( .A(n1602), .B(n1448), .Y(n1463) );
  AOI21X1 U1965 ( .A(n2304), .B(n1742), .C(n1942), .Y(n2302) );
  NAND3X1 U1966 ( .A(n1847), .B(n2305), .C(n1849), .Y(n1742) );
  NAND3X1 U1967 ( .A(n1378), .B(n1939), .C(n2306), .Y(n2304) );
  AOI21X1 U1968 ( .A(n2307), .B(n2308), .C(n2309), .Y(n2306) );
  INVX1 U1969 ( .A(n1585), .Y(n2309) );
  NAND3X1 U1970 ( .A(n2022), .B(n1633), .C(n1945), .Y(n1585) );
  OAI21X1 U1971 ( .A(n2162), .B(n2310), .C(n2311), .Y(n2308) );
  AND2X1 U1972 ( .A(n1640), .B(n1390), .Y(n2311) );
  NAND2X1 U1973 ( .A(n1526), .B(n2029), .Y(n1640) );
  AOI21X1 U1974 ( .A(n2034), .B(n2312), .C(n2313), .Y(n2310) );
  INVX1 U1975 ( .A(n1393), .Y(n2313) );
  NAND3X1 U1976 ( .A(n2287), .B(n1982), .C(n1679), .Y(n1393) );
  OAI21X1 U1977 ( .A(n2314), .B(n2315), .C(n2316), .Y(n2312) );
  INVX1 U1978 ( .A(n1592), .Y(n2316) );
  NAND2X1 U1979 ( .A(n1394), .B(n1806), .Y(n1592) );
  AND2X1 U1980 ( .A(n2209), .B(n1760), .Y(n1394) );
  NAND3X1 U1981 ( .A(n2287), .B(n2235), .C(n2317), .Y(n1760) );
  NOR2X1 U1982 ( .A(n1451), .B(n2237), .Y(n2317) );
  NAND2X1 U1983 ( .A(n2170), .B(n1591), .Y(n2315) );
  NAND3X1 U1984 ( .A(n1923), .B(n1250), .C(n1847), .Y(n2170) );
  AOI21X1 U1985 ( .A(n1398), .B(n2318), .C(n1597), .Y(n2314) );
  OAI21X1 U1986 ( .A(n2319), .B(n2320), .C(n1758), .Y(n2318) );
  INVX1 U1987 ( .A(n1907), .Y(n1758) );
  NAND2X1 U1988 ( .A(n2065), .B(n1404), .Y(n1907) );
  NAND3X1 U1989 ( .A(n1938), .B(n1987), .C(n1986), .Y(n1404) );
  INVX1 U1990 ( .A(n1459), .Y(n2320) );
  AOI21X1 U1991 ( .A(n2176), .B(n2321), .C(n1763), .Y(n2319) );
  INVX1 U1992 ( .A(n1914), .Y(n1763) );
  NAND3X1 U1993 ( .A(n1986), .B(n1457), .C(n1924), .Y(n1914) );
  OAI21X1 U1994 ( .A(n2322), .B(n2323), .C(n2324), .Y(n2321) );
  NOR2X1 U1995 ( .A(n2064), .B(n2048), .Y(n2324) );
  NOR2X1 U1996 ( .A(n1937), .B(n2208), .Y(n2048) );
  AOI21X1 U1997 ( .A(n1799), .B(n1751), .C(n1937), .Y(n2064) );
  NAND2X1 U1998 ( .A(n1615), .B(n1410), .Y(n2323) );
  AOI21X1 U1999 ( .A(n2325), .B(n1419), .C(n2326), .Y(n2322) );
  NAND2X1 U2000 ( .A(n1611), .B(n2187), .Y(n2326) );
  NAND2X1 U2001 ( .A(n2290), .B(n1964), .Y(n1419) );
  OAI21X1 U2002 ( .A(n1638), .B(n2327), .C(n2328), .Y(n2325) );
  INVX1 U2003 ( .A(n1617), .Y(n2328) );
  NAND2X1 U2004 ( .A(n1421), .B(n1773), .Y(n1617) );
  NAND3X1 U2005 ( .A(n1447), .B(n1982), .C(n1526), .Y(n1773) );
  OAI21X1 U2006 ( .A(n2329), .B(n2330), .C(n1778), .Y(n2327) );
  INVX1 U2007 ( .A(n1926), .Y(n2330) );
  NAND3X1 U2008 ( .A(n2260), .B(n1982), .C(n1526), .Y(n1926) );
  AND2X1 U2009 ( .A(n2331), .B(n1780), .Y(n2329) );
  OAI21X1 U2010 ( .A(n1795), .B(n2332), .C(n1932), .Y(n2331) );
  AOI21X1 U2011 ( .A(n2333), .B(n2334), .C(n2202), .Y(n2332) );
  INVX1 U2012 ( .A(n1441), .Y(n2202) );
  NAND3X1 U2013 ( .A(n1829), .B(n1986), .C(n1632), .Y(n1441) );
  OAI21X1 U2014 ( .A(n2335), .B(n2336), .C(n2337), .Y(n2334) );
  NOR2X1 U2015 ( .A(state[4]), .B(n1797), .Y(n2337) );
  INVX1 U2016 ( .A(n2060), .Y(n1797) );
  NAND2X1 U2017 ( .A(n1630), .B(n2338), .Y(n2336) );
  NAND3X1 U2018 ( .A(next_byte[6]), .B(n2339), .C(n2340), .Y(n2335) );
  NAND2X1 U2019 ( .A(n2052), .B(n2191), .Y(n1638) );
  NAND3X1 U2020 ( .A(n1993), .B(n1986), .C(n1454), .Y(n2191) );
  NOR2X1 U2021 ( .A(n2341), .B(n2342), .Y(n1454) );
  NOR2X1 U2022 ( .A(n1582), .B(n1893), .Y(n2307) );
  INVX1 U2023 ( .A(n1386), .Y(n1582) );
  NAND3X1 U2024 ( .A(n2118), .B(n1601), .C(n1768), .Y(n1386) );
  NAND3X1 U2025 ( .A(n1982), .B(n1416), .C(n1945), .Y(n1378) );
  NAND2X1 U2026 ( .A(n2211), .B(n2068), .Y(n2297) );
  NAND2X1 U2027 ( .A(n2021), .B(n1251), .Y(n2068) );
  NAND3X1 U2028 ( .A(n1964), .B(n1414), .C(n1941), .Y(n2211) );
  INVX1 U2029 ( .A(n1730), .Y(n1879) );
  NAND3X1 U2030 ( .A(n1922), .B(n1929), .C(n1849), .Y(n1730) );
  AND2X1 U2031 ( .A(n1467), .B(n1723), .Y(n2294) );
  NAND2X1 U2032 ( .A(n2343), .B(n1650), .Y(n1723) );
  NAND2X1 U2033 ( .A(n2344), .B(n1355), .Y(n1546) );
  NAND2X1 U2034 ( .A(n1455), .B(n2290), .Y(n1355) );
  NAND3X1 U2035 ( .A(n1602), .B(n1633), .C(n2218), .Y(n1543) );
  INVX1 U2036 ( .A(n1541), .Y(n2000) );
  NAND3X1 U2037 ( .A(n1829), .B(n1982), .C(n2345), .Y(n1541) );
  AND2X1 U2038 ( .A(n1538), .B(n2215), .Y(n2275) );
  NAND3X1 U2039 ( .A(n2345), .B(n2227), .C(n2346), .Y(n2215) );
  NOR2X1 U2040 ( .A(state[1]), .B(n1637), .Y(n2346) );
  INVX1 U2041 ( .A(n2347), .Y(n2345) );
  NAND3X1 U2042 ( .A(n2348), .B(next_byte[3]), .C(n2349), .Y(n2347) );
  NOR2X1 U2043 ( .A(n2350), .B(n2351), .Y(n2349) );
  NOR2X1 U2044 ( .A(next_byte[6]), .B(n2339), .Y(n2348) );
  INVX1 U2045 ( .A(n1328), .Y(n2273) );
  NAND3X1 U2046 ( .A(n1704), .B(n1632), .C(n2352), .Y(n1328) );
  NOR2X1 U2047 ( .A(n1451), .B(n2256), .Y(n2352) );
  INVX1 U2048 ( .A(n2115), .Y(n2268) );
  NOR2X1 U2049 ( .A(n1751), .B(n2111), .Y(n2266) );
  INVX1 U2050 ( .A(n2353), .Y(n2075) );
  NOR2X1 U2051 ( .A(n1683), .B(n2100), .Y(n2253) );
  INVX1 U2052 ( .A(n1837), .Y(n2100) );
  INVX1 U2053 ( .A(n1305), .Y(n1683) );
  NAND2X1 U2054 ( .A(n2354), .B(n2355), .Y(n1305) );
  INVX1 U2055 ( .A(n1302), .Y(n1682) );
  NAND3X1 U2056 ( .A(n1705), .B(n2057), .C(n2106), .Y(n1302) );
  INVX1 U2057 ( .A(n1276), .Y(n2242) );
  AND2X1 U2058 ( .A(n1650), .B(n1944), .Y(n2238) );
  INVX1 U2059 ( .A(n1663), .Y(n1272) );
  NAND2X1 U2060 ( .A(n2290), .B(n1650), .Y(n1663) );
  AND2X1 U2061 ( .A(n1250), .B(n1678), .Y(n2290) );
  INVX1 U2062 ( .A(n1956), .Y(n2231) );
  NAND3X1 U2063 ( .A(n2085), .B(n1678), .C(n1768), .Y(n1956) );
  NOR2X1 U2064 ( .A(n1264), .B(n2076), .Y(n2228) );
  INVX1 U2065 ( .A(n1480), .Y(n1264) );
  NAND3X1 U2066 ( .A(n1650), .B(n2356), .C(n1250), .Y(n1480) );
  NAND3X1 U2067 ( .A(n2357), .B(n1647), .C(n2358), .Y(n1234) );
  MUX2X1 U2068 ( .B(n1263), .A(state[2]), .S(n1259), .Y(n2358) );
  INVX1 U2069 ( .A(n1479), .Y(n1263) );
  NAND3X1 U2070 ( .A(n2250), .B(n1678), .C(n1804), .Y(n1479) );
  NAND3X1 U2071 ( .A(n2072), .B(n1677), .C(n2359), .Y(n1647) );
  NOR2X1 U2072 ( .A(n1259), .B(n2360), .Y(n2359) );
  INVX1 U2073 ( .A(en), .Y(n1259) );
  NOR2X1 U2074 ( .A(n1636), .B(n2361), .Y(n1677) );
  NAND3X1 U2075 ( .A(n2362), .B(n1952), .C(n2363), .Y(n2357) );
  INVX1 U2076 ( .A(n1955), .Y(n2363) );
  NAND2X1 U2077 ( .A(en), .B(n1652), .Y(n1955) );
  NAND3X1 U2078 ( .A(n2213), .B(n2364), .C(n2272), .Y(n1652) );
  NAND2X1 U2079 ( .A(n2213), .B(n2343), .Y(n1952) );
  OAI21X1 U2080 ( .A(n2365), .B(n2076), .C(n1815), .Y(n2362) );
  NAND3X1 U2081 ( .A(n1986), .B(n2272), .C(n2043), .Y(n1815) );
  INVX1 U2082 ( .A(n1266), .Y(n2076) );
  NAND3X1 U2083 ( .A(n1929), .B(n2355), .C(n1796), .Y(n1266) );
  AOI21X1 U2084 ( .A(n1654), .B(n2366), .C(n2367), .Y(n2365) );
  INVX1 U2085 ( .A(n1270), .Y(n2367) );
  NAND2X1 U2086 ( .A(n2354), .B(n2106), .Y(n1270) );
  OAI21X1 U2087 ( .A(n1961), .B(n2368), .C(n2369), .Y(n2366) );
  AND2X1 U2088 ( .A(n1474), .B(n2086), .Y(n2369) );
  NAND3X1 U2089 ( .A(n1633), .B(n1501), .C(n2085), .Y(n2086) );
  NAND3X1 U2090 ( .A(n2089), .B(n1414), .C(n1416), .Y(n1474) );
  NAND2X1 U2091 ( .A(n2370), .B(n1471), .Y(n2368) );
  NAND3X1 U2092 ( .A(n1982), .B(n1629), .C(n2204), .Y(n1471) );
  OAI21X1 U2093 ( .A(n1276), .B(n2371), .C(n1665), .Y(n2370) );
  NOR2X1 U2094 ( .A(n1490), .B(n2244), .Y(n1665) );
  INVX1 U2095 ( .A(n1824), .Y(n2244) );
  NAND3X1 U2096 ( .A(n2089), .B(n2085), .C(n1982), .Y(n1824) );
  INVX1 U2097 ( .A(n1472), .Y(n1490) );
  NAND3X1 U2098 ( .A(n1944), .B(n1982), .C(n1457), .Y(n1472) );
  NOR2X1 U2099 ( .A(n2342), .B(n2361), .Y(n1944) );
  OAI21X1 U2100 ( .A(n2372), .B(n1496), .C(n1668), .Y(n2371) );
  NAND2X1 U2101 ( .A(n1829), .B(n1813), .Y(n1668) );
  INVX1 U2102 ( .A(n2247), .Y(n1496) );
  NAND3X1 U2103 ( .A(n1804), .B(n2250), .C(n1982), .Y(n2247) );
  AOI21X1 U2104 ( .A(n1669), .B(n2373), .C(n2374), .Y(n2372) );
  INVX1 U2105 ( .A(n1283), .Y(n2374) );
  NAND3X1 U2106 ( .A(n2272), .B(n1982), .C(n2158), .Y(n1283) );
  OAI21X1 U2107 ( .A(n1675), .B(n2375), .C(n1289), .Y(n2373) );
  NAND3X1 U2108 ( .A(n1829), .B(n2376), .C(n2377), .Y(n1289) );
  NOR2X1 U2109 ( .A(n2341), .B(n1637), .Y(n2377) );
  AOI21X1 U2110 ( .A(n2378), .B(n1298), .C(n1830), .Y(n2375) );
  INVX1 U2111 ( .A(n1504), .Y(n1830) );
  NAND3X1 U2112 ( .A(n2069), .B(state[2]), .C(n2354), .Y(n1504) );
  NAND3X1 U2113 ( .A(n2227), .B(n1796), .C(n2379), .Y(n1298) );
  NOR2X1 U2114 ( .A(n1451), .B(n1476), .Y(n2379) );
  OAI21X1 U2115 ( .A(n1974), .B(n2380), .C(n1971), .Y(n2378) );
  NAND2X1 U2116 ( .A(n1447), .B(n1500), .Y(n1971) );
  NAND2X1 U2117 ( .A(n2381), .B(n1837), .Y(n2380) );
  NAND3X1 U2118 ( .A(n2022), .B(n2070), .C(n1922), .Y(n1837) );
  NAND3X1 U2119 ( .A(n2353), .B(n1681), .C(n2382), .Y(n2381) );
  OAI21X1 U2120 ( .A(n2383), .B(n1839), .C(n1514), .Y(n2382) );
  NAND3X1 U2121 ( .A(n1704), .B(n1629), .C(n2210), .Y(n1514) );
  INVX1 U2122 ( .A(n1306), .Y(n1839) );
  NAND3X1 U2123 ( .A(n1601), .B(n1250), .C(n1940), .Y(n1306) );
  AOI21X1 U2124 ( .A(n1842), .B(n2384), .C(n1978), .Y(n2383) );
  INVX1 U2125 ( .A(n1313), .Y(n1978) );
  NAND3X1 U2126 ( .A(n2250), .B(n1629), .C(n1601), .Y(n1313) );
  NAND3X1 U2127 ( .A(n1980), .B(n1643), .C(n2385), .Y(n2384) );
  OAI21X1 U2128 ( .A(n2110), .B(n2111), .C(n2386), .Y(n2385) );
  AOI21X1 U2129 ( .A(n2387), .B(n2115), .C(n1519), .Y(n2386) );
  INVX1 U2130 ( .A(n2388), .Y(n1519) );
  NAND3X1 U2131 ( .A(n1964), .B(n1987), .C(n1986), .Y(n2388) );
  NAND3X1 U2132 ( .A(n1982), .B(n1250), .C(n2389), .Y(n2115) );
  OAI21X1 U2133 ( .A(n1326), .B(n2390), .C(n1325), .Y(n2387) );
  NAND3X1 U2134 ( .A(n1986), .B(n2085), .C(n2158), .Y(n1325) );
  AOI21X1 U2135 ( .A(n2391), .B(n1333), .C(n1531), .Y(n2390) );
  INVX1 U2136 ( .A(n1330), .Y(n1531) );
  NAND3X1 U2137 ( .A(n2069), .B(n1250), .C(n1923), .Y(n1330) );
  NAND3X1 U2138 ( .A(n1796), .B(n1601), .C(n2089), .Y(n1333) );
  OAI21X1 U2139 ( .A(n2392), .B(n2393), .C(n1538), .Y(n2391) );
  NAND3X1 U2140 ( .A(n2112), .B(n1633), .C(n2354), .Y(n1538) );
  AOI21X1 U2141 ( .A(n1943), .B(n2394), .C(n2125), .Y(n2393) );
  INVX1 U2142 ( .A(n1337), .Y(n2125) );
  NAND3X1 U2143 ( .A(n1923), .B(n2072), .C(n2127), .Y(n1337) );
  INVX1 U2144 ( .A(n2395), .Y(n1923) );
  NAND3X1 U2145 ( .A(n2396), .B(n1544), .C(n1714), .Y(n2394) );
  NOR2X1 U2146 ( .A(n2282), .B(n1339), .Y(n1714) );
  INVX1 U2147 ( .A(n1861), .Y(n1339) );
  NAND3X1 U2148 ( .A(n2272), .B(n1601), .C(n2158), .Y(n1861) );
  INVX1 U2149 ( .A(n1347), .Y(n2282) );
  NAND3X1 U2150 ( .A(n1986), .B(n1629), .C(n1768), .Y(n1347) );
  NAND2X1 U2151 ( .A(n1768), .B(n1963), .Y(n1544) );
  OAI21X1 U2152 ( .A(n2397), .B(n1720), .C(n2398), .Y(n2396) );
  AND2X1 U2153 ( .A(n1343), .B(n2004), .Y(n2398) );
  NAND3X1 U2154 ( .A(n2066), .B(n2022), .C(n1706), .Y(n2004) );
  NAND3X1 U2155 ( .A(n2118), .B(n1929), .C(n1706), .Y(n1343) );
  INVX1 U2156 ( .A(n2344), .Y(n1720) );
  NAND3X1 U2157 ( .A(n1633), .B(n2213), .C(n2022), .Y(n2344) );
  AOI21X1 U2158 ( .A(n1551), .B(n2399), .C(n2400), .Y(n2397) );
  INVX1 U2159 ( .A(n1349), .Y(n2400) );
  NAND3X1 U2160 ( .A(n1601), .B(n1629), .C(n1457), .Y(n1349) );
  OAI21X1 U2161 ( .A(n2401), .B(n2402), .C(n1867), .Y(n2399) );
  NOR2X1 U2162 ( .A(n2403), .B(n2292), .Y(n1867) );
  INVX1 U2163 ( .A(n2404), .Y(n2292) );
  NAND3X1 U2164 ( .A(n1982), .B(n1650), .C(n1526), .Y(n2404) );
  INVX1 U2165 ( .A(n1357), .Y(n2403) );
  NAND3X1 U2166 ( .A(n1650), .B(n1414), .C(n1628), .Y(n1357) );
  NAND2X1 U2167 ( .A(n1873), .B(n1468), .Y(n2402) );
  NAND3X1 U2168 ( .A(n1250), .B(n1414), .C(n1993), .Y(n1468) );
  NAND3X1 U2169 ( .A(n1804), .B(n1415), .C(n1601), .Y(n1873) );
  AOI21X1 U2170 ( .A(n1728), .B(n2405), .C(n1870), .Y(n2401) );
  INVX1 U2171 ( .A(n2137), .Y(n1870) );
  NAND2X1 U2172 ( .A(n2343), .B(n1501), .Y(n2137) );
  NOR2X1 U2173 ( .A(n2180), .B(n2120), .Y(n1501) );
  NOR2X1 U2174 ( .A(n2171), .B(n2406), .Y(n2343) );
  INVX1 U2175 ( .A(n1803), .Y(n2171) );
  NOR2X1 U2176 ( .A(n1636), .B(n2407), .Y(n1803) );
  OAI21X1 U2177 ( .A(n2408), .B(n2409), .C(n2212), .Y(n2405) );
  NAND3X1 U2178 ( .A(n2106), .B(n2305), .C(n2410), .Y(n2212) );
  NOR2X1 U2179 ( .A(n2411), .B(n1790), .Y(n2410) );
  AND2X1 U2180 ( .A(n1922), .B(n2116), .Y(n2106) );
  NAND2X1 U2181 ( .A(n1467), .B(n1466), .Y(n2409) );
  NAND3X1 U2182 ( .A(n2056), .B(n2085), .C(n1704), .Y(n1466) );
  NAND3X1 U2183 ( .A(n1704), .B(n2056), .C(n2412), .Y(n1467) );
  NOR2X1 U2184 ( .A(n1636), .B(n1790), .Y(n2412) );
  NAND3X1 U2185 ( .A(next_byte[3]), .B(n2413), .C(next_byte[4]), .Y(n1636) );
  AOI21X1 U2186 ( .A(n1368), .B(n2414), .C(n2016), .Y(n2408) );
  INVX1 U2187 ( .A(n1556), .Y(n2016) );
  NAND3X1 U2188 ( .A(n1601), .B(n1250), .C(n1455), .Y(n1556) );
  OAI21X1 U2189 ( .A(n1881), .B(n2415), .C(n1369), .Y(n2414) );
  NAND3X1 U2190 ( .A(n1796), .B(n2057), .C(n1706), .Y(n1369) );
  NOR2X1 U2191 ( .A(n2416), .B(state[2]), .Y(n1706) );
  OAI21X1 U2192 ( .A(n2417), .B(n2418), .C(n2145), .Y(n2415) );
  NAND3X1 U2193 ( .A(n1922), .B(n1629), .C(n2073), .Y(n2145) );
  NAND2X1 U2194 ( .A(n1740), .B(n2020), .Y(n2418) );
  NAND3X1 U2195 ( .A(n1633), .B(n1796), .C(n2389), .Y(n2020) );
  NAND3X1 U2196 ( .A(n1895), .B(n1633), .C(n2260), .Y(n1740) );
  AOI21X1 U2197 ( .A(n2419), .B(n2420), .C(n1641), .Y(n2417) );
  INVX1 U2198 ( .A(n1464), .Y(n1641) );
  NAND3X1 U2199 ( .A(n2204), .B(n1414), .C(n1924), .Y(n1464) );
  OAI21X1 U2200 ( .A(n2421), .B(n1385), .C(n2028), .Y(n2420) );
  AND2X1 U2201 ( .A(n1574), .B(n1939), .Y(n2028) );
  NAND2X1 U2202 ( .A(n1940), .B(n1448), .Y(n1939) );
  NOR2X1 U2203 ( .A(n1751), .B(n1451), .Y(n1448) );
  NAND2X1 U2204 ( .A(n2155), .B(n1813), .Y(n1574) );
  NOR2X1 U2205 ( .A(n2208), .B(n1451), .Y(n1813) );
  AND2X1 U2206 ( .A(n2248), .B(n1457), .Y(n1385) );
  NOR2X1 U2207 ( .A(n1799), .B(n1254), .Y(n2248) );
  AOI21X1 U2208 ( .A(n1898), .B(n2422), .C(n1893), .Y(n2421) );
  INVX1 U2209 ( .A(n1588), .Y(n1893) );
  NAND3X1 U2210 ( .A(n1705), .B(n2069), .C(n2073), .Y(n1588) );
  NAND3X1 U2211 ( .A(n1390), .B(n1461), .C(n2423), .Y(n2422) );
  OAI21X1 U2212 ( .A(n2162), .B(n2424), .C(n1589), .Y(n2423) );
  NAND2X1 U2213 ( .A(n1988), .B(n1963), .Y(n1589) );
  INVX1 U2214 ( .A(n2425), .Y(n2424) );
  OAI21X1 U2215 ( .A(n2426), .B(n2427), .C(n1902), .Y(n2425) );
  AND2X1 U2216 ( .A(n2034), .B(n1806), .Y(n1902) );
  NAND2X1 U2217 ( .A(n1963), .B(n1650), .Y(n1806) );
  NOR2X1 U2218 ( .A(n2428), .B(state[1]), .Y(n1650) );
  NAND3X1 U2219 ( .A(n2178), .B(n2070), .C(n2429), .Y(n2034) );
  NOR2X1 U2220 ( .A(n2416), .B(n2205), .Y(n2429) );
  INVX1 U2221 ( .A(n2430), .Y(n2205) );
  INVX1 U2222 ( .A(n2360), .Y(n2070) );
  INVX1 U2223 ( .A(n2341), .Y(n2178) );
  OAI21X1 U2224 ( .A(n2431), .B(n1597), .C(n2035), .Y(n2427) );
  NOR2X1 U2225 ( .A(n1755), .B(n1392), .Y(n2035) );
  INVX1 U2226 ( .A(n2432), .Y(n1392) );
  NAND3X1 U2227 ( .A(n2030), .B(n2305), .C(n1930), .Y(n2432) );
  NOR2X1 U2228 ( .A(n2433), .B(n1476), .Y(n1922) );
  INVX1 U2229 ( .A(n1591), .Y(n1755) );
  NAND3X1 U2230 ( .A(n1993), .B(n1678), .C(n1628), .Y(n1591) );
  INVX1 U2231 ( .A(n1909), .Y(n1597) );
  NAND3X1 U2232 ( .A(n2272), .B(n1982), .C(n1602), .Y(n1909) );
  AOI21X1 U2233 ( .A(n2434), .B(n1401), .C(n2435), .Y(n2431) );
  INVX1 U2234 ( .A(n1398), .Y(n2435) );
  NAND3X1 U2235 ( .A(n1416), .B(n1678), .C(n1938), .Y(n1398) );
  NOR2X1 U2236 ( .A(n2436), .B(n2341), .Y(n1416) );
  NAND3X1 U2237 ( .A(n2272), .B(n1601), .C(n2260), .Y(n1401) );
  AND2X1 U2238 ( .A(n2066), .B(n1814), .Y(n2260) );
  OAI21X1 U2239 ( .A(n2437), .B(n2438), .C(n2065), .Y(n2434) );
  NAND3X1 U2240 ( .A(n1847), .B(n2272), .C(n2073), .Y(n2065) );
  INVX1 U2241 ( .A(n2439), .Y(n2073) );
  NAND2X1 U2242 ( .A(n1802), .B(n1459), .Y(n2438) );
  NAND3X1 U2243 ( .A(n2227), .B(n2072), .C(n2287), .Y(n1459) );
  NAND2X1 U2244 ( .A(n1805), .B(n2022), .Y(n1802) );
  NOR2X1 U2245 ( .A(n1789), .B(n2440), .Y(n1805) );
  AOI21X1 U2246 ( .A(n1918), .B(n2441), .C(n1765), .Y(n2437) );
  OAI21X1 U2247 ( .A(n1751), .B(n1937), .C(n2176), .Y(n1765) );
  NAND3X1 U2248 ( .A(n2356), .B(n1415), .C(n1924), .Y(n2176) );
  NAND2X1 U2249 ( .A(n1986), .B(n1415), .Y(n1937) );
  OAI21X1 U2250 ( .A(n2207), .B(n2442), .C(n2443), .Y(n2441) );
  NOR2X1 U2251 ( .A(n2045), .B(n1408), .Y(n2443) );
  INVX1 U2252 ( .A(n1611), .Y(n1408) );
  NAND3X1 U2253 ( .A(n1705), .B(n1982), .C(n1940), .Y(n1611) );
  NOR2X1 U2254 ( .A(n2395), .B(n1476), .Y(n1940) );
  INVX1 U2255 ( .A(n1406), .Y(n2045) );
  NAND3X1 U2256 ( .A(n1679), .B(n1453), .C(n2444), .Y(n1406) );
  NOR2X1 U2257 ( .A(n2445), .B(n1451), .Y(n2444) );
  INVX1 U2258 ( .A(n2446), .Y(n1453) );
  AOI21X1 U2259 ( .A(n2447), .B(n1420), .C(n2448), .Y(n2442) );
  INVX1 U2260 ( .A(n2187), .Y(n2448) );
  NAND3X1 U2261 ( .A(n1804), .B(n1415), .C(n1633), .Y(n2187) );
  NAND3X1 U2262 ( .A(n2043), .B(n1601), .C(n2030), .Y(n1420) );
  OAI21X1 U2263 ( .A(n2053), .B(n2449), .C(n2206), .Y(n2447) );
  NAND3X1 U2264 ( .A(n2356), .B(n1804), .C(n2213), .Y(n2206) );
  AOI21X1 U2265 ( .A(n2450), .B(n1778), .C(n2451), .Y(n2449) );
  INVX1 U2266 ( .A(n2052), .Y(n2451) );
  NAND3X1 U2267 ( .A(n2056), .B(n1929), .C(n1924), .Y(n2052) );
  NAND3X1 U2268 ( .A(n1988), .B(n1601), .C(n1994), .Y(n1778) );
  NOR2X1 U2269 ( .A(n2361), .B(n2411), .Y(n1994) );
  NOR2X1 U2270 ( .A(n2428), .B(n1476), .Y(n1988) );
  OAI21X1 U2271 ( .A(n2452), .B(n1783), .C(n1780), .Y(n2450) );
  NAND3X1 U2272 ( .A(n1829), .B(n1678), .C(n1628), .Y(n1780) );
  NOR2X1 U2273 ( .A(n2256), .B(n2104), .Y(n1829) );
  NAND2X1 U2274 ( .A(n1932), .B(n1433), .Y(n1783) );
  NAND3X1 U2275 ( .A(n1986), .B(n2089), .C(n1632), .Y(n1433) );
  NOR2X1 U2276 ( .A(n1790), .B(n2445), .Y(n1632) );
  NAND3X1 U2277 ( .A(n1986), .B(n2453), .C(n2454), .Y(n1932) );
  NOR2X1 U2278 ( .A(n2361), .B(n1659), .Y(n2454) );
  AOI21X1 U2279 ( .A(n2333), .B(n2455), .C(n1795), .Y(n2452) );
  INVX1 U2280 ( .A(n1436), .Y(n1795) );
  NAND3X1 U2281 ( .A(n2364), .B(n1415), .C(n1924), .Y(n1436) );
  NOR2X1 U2282 ( .A(n2446), .B(n2436), .Y(n1924) );
  INVX1 U2283 ( .A(n1253), .Y(n1415) );
  OAI21X1 U2284 ( .A(state[2]), .B(n1631), .C(n2060), .Y(n2455) );
  NAND3X1 U2285 ( .A(n1630), .B(n2456), .C(n2430), .Y(n2060) );
  INVX1 U2286 ( .A(n2457), .Y(n1630) );
  INVX1 U2287 ( .A(n1446), .Y(n1631) );
  NAND3X1 U2288 ( .A(n1457), .B(n1633), .C(n2030), .Y(n1446) );
  NOR2X1 U2289 ( .A(n1476), .B(n2360), .Y(n1457) );
  INVX1 U2290 ( .A(n1439), .Y(n2333) );
  OAI21X1 U2291 ( .A(n1799), .B(n2457), .C(n2203), .Y(n1439) );
  NAND3X1 U2292 ( .A(n2287), .B(n1601), .C(n2389), .Y(n2203) );
  AND2X1 U2293 ( .A(n2338), .B(n2453), .Y(n2287) );
  INVX1 U2294 ( .A(n2436), .Y(n2453) );
  NAND2X1 U2295 ( .A(n1768), .B(n1414), .Y(n2457) );
  NOR2X1 U2296 ( .A(n2439), .B(n1476), .Y(n1768) );
  INVX1 U2297 ( .A(n1421), .Y(n2053) );
  NAND3X1 U2298 ( .A(n2458), .B(n2456), .C(n2459), .Y(n1421) );
  AND2X1 U2299 ( .A(n1982), .B(n2043), .Y(n2459) );
  NOR2X1 U2300 ( .A(n2104), .B(n2180), .Y(n2043) );
  INVX1 U2301 ( .A(n2221), .Y(n2180) );
  NOR2X1 U2302 ( .A(state[1]), .B(state[2]), .Y(n2221) );
  INVX1 U2303 ( .A(n2361), .Y(n2456) );
  INVX1 U2304 ( .A(n1615), .Y(n2207) );
  NAND3X1 U2305 ( .A(n2072), .B(n2057), .C(n1849), .Y(n1615) );
  AND2X1 U2306 ( .A(n1250), .B(n2116), .Y(n1849) );
  NOR2X1 U2307 ( .A(n1612), .B(n2460), .Y(n1918) );
  INVX1 U2308 ( .A(n1771), .Y(n2460) );
  NAND2X1 U2309 ( .A(n1455), .B(n1500), .Y(n1771) );
  INVX1 U2310 ( .A(n1286), .Y(n1500) );
  NAND2X1 U2311 ( .A(n1986), .B(n1250), .Y(n1286) );
  INVX1 U2312 ( .A(n1410), .Y(n1612) );
  NAND3X1 U2313 ( .A(n2210), .B(n2057), .C(n1526), .Y(n1410) );
  NOR2X1 U2314 ( .A(n2195), .B(state[2]), .Y(n2210) );
  INVX1 U2315 ( .A(n2069), .Y(n2195) );
  NAND2X1 U2316 ( .A(n1595), .B(n2209), .Y(n2426) );
  NAND3X1 U2317 ( .A(n2085), .B(n1414), .C(n1938), .Y(n2209) );
  NAND3X1 U2318 ( .A(n2430), .B(n1938), .C(n2197), .Y(n1595) );
  NOR2X1 U2319 ( .A(n2407), .B(n1451), .Y(n2197) );
  NOR2X1 U2320 ( .A(n2461), .B(next_byte[4]), .Y(n2430) );
  INVX1 U2321 ( .A(n1639), .Y(n2162) );
  NAND3X1 U2322 ( .A(n2158), .B(n1678), .C(n2030), .Y(n1639) );
  AND2X1 U2323 ( .A(n2338), .B(n2376), .Y(n2030) );
  INVX1 U2324 ( .A(n2342), .Y(n2376) );
  OR2X1 U2325 ( .A(n1752), .B(n2110), .Y(n1461) );
  INVX1 U2326 ( .A(n2029), .Y(n1752) );
  NOR2X1 U2327 ( .A(n2440), .B(n2462), .Y(n2029) );
  NAND3X1 U2328 ( .A(n2213), .B(n1414), .C(n1796), .Y(n1390) );
  NOR2X1 U2329 ( .A(n2341), .B(n2411), .Y(n1796) );
  NAND3X1 U2330 ( .A(n2463), .B(n2464), .C(n2465), .Y(n2341) );
  INVX1 U2331 ( .A(n2462), .Y(n2213) );
  NAND3X1 U2332 ( .A(n2466), .B(n2467), .C(state[2]), .Y(n2462) );
  NAND3X1 U2333 ( .A(n2089), .B(n2356), .C(n1526), .Y(n1898) );
  AND2X1 U2334 ( .A(n1570), .B(n2153), .Y(n2419) );
  INVX1 U2335 ( .A(n1942), .Y(n2153) );
  NOR2X1 U2336 ( .A(n2468), .B(n2230), .Y(n1942) );
  INVX1 U2337 ( .A(n2156), .Y(n2230) );
  NAND2X1 U2338 ( .A(n1602), .B(n2113), .Y(n1570) );
  AND2X1 U2339 ( .A(n1987), .B(n1414), .Y(n2113) );
  OAI21X1 U2340 ( .A(n1565), .B(n1566), .C(n2019), .Y(n1881) );
  NAND2X1 U2341 ( .A(n2021), .B(n1804), .Y(n2019) );
  INVX1 U2342 ( .A(n2208), .Y(n1804) );
  NAND3X1 U2343 ( .A(n2469), .B(n2458), .C(next_byte[1]), .Y(n2208) );
  NOR2X1 U2344 ( .A(n1800), .B(n1253), .Y(n2021) );
  NAND3X1 U2345 ( .A(state[2]), .B(n2466), .C(state[3]), .Y(n1253) );
  INVX1 U2346 ( .A(n2354), .Y(n1566) );
  NOR2X1 U2347 ( .A(n2237), .B(n1799), .Y(n2354) );
  INVX1 U2348 ( .A(n2056), .Y(n1565) );
  NAND3X1 U2349 ( .A(n1704), .B(n2355), .C(n1628), .Y(n1368) );
  AND2X1 U2350 ( .A(n2338), .B(n1456), .Y(n1628) );
  NAND3X1 U2351 ( .A(n2355), .B(n2057), .C(n2272), .Y(n1728) );
  NAND3X1 U2352 ( .A(n2204), .B(n1633), .C(n1941), .Y(n1551) );
  NOR2X1 U2353 ( .A(n2411), .B(n2407), .Y(n1941) );
  NOR2X1 U2354 ( .A(n2129), .B(n1539), .Y(n1943) );
  INVX1 U2355 ( .A(n2470), .Y(n1539) );
  NAND3X1 U2356 ( .A(n1895), .B(n1986), .C(n1602), .Y(n2470) );
  NAND3X1 U2357 ( .A(state[0]), .B(n2225), .C(state[6]), .Y(n2440) );
  INVX1 U2358 ( .A(n1998), .Y(n2129) );
  NAND3X1 U2359 ( .A(n2089), .B(n2364), .C(n1895), .Y(n1998) );
  AND2X1 U2360 ( .A(n2338), .B(n2458), .Y(n1895) );
  INVX1 U2361 ( .A(n2411), .Y(n2458) );
  AND2X1 U2362 ( .A(n2469), .B(n2463), .Y(n2338) );
  INVX1 U2363 ( .A(n1659), .Y(n2089) );
  NAND3X1 U2364 ( .A(n2116), .B(n2467), .C(n2466), .Y(n1659) );
  INVX1 U2365 ( .A(n1535), .Y(n2392) );
  NAND3X1 U2366 ( .A(n2127), .B(n2356), .C(n1602), .Y(n1535) );
  INVX1 U2367 ( .A(n2433), .Y(n2356) );
  INVX1 U2368 ( .A(n2471), .Y(n2127) );
  INVX1 U2369 ( .A(n2472), .Y(n1326) );
  NAND3X1 U2370 ( .A(n1633), .B(n2250), .C(n2272), .Y(n2472) );
  AND2X1 U2371 ( .A(n1814), .B(n2057), .Y(n2250) );
  NAND2X1 U2372 ( .A(n1447), .B(n1601), .Y(n2111) );
  NOR2X1 U2373 ( .A(n1526), .B(n2022), .Y(n2110) );
  NOR2X1 U2374 ( .A(n2436), .B(n2407), .Y(n1526) );
  NAND3X1 U2375 ( .A(next_byte[5]), .B(n2473), .C(n2340), .Y(n2436) );
  NAND3X1 U2376 ( .A(n1987), .B(n1678), .C(n2389), .Y(n1643) );
  INVX1 U2377 ( .A(n1789), .Y(n2389) );
  NAND2X1 U2378 ( .A(n1929), .B(n1814), .Y(n1789) );
  NAND3X1 U2379 ( .A(n1250), .B(n2364), .C(n1602), .Y(n1980) );
  INVX1 U2380 ( .A(n2468), .Y(n1602) );
  NAND3X1 U2381 ( .A(n2466), .B(n2116), .C(state[3]), .Y(n2468) );
  AND2X1 U2382 ( .A(n2474), .B(n1476), .Y(n2466) );
  INVX1 U2383 ( .A(n1807), .Y(n2364) );
  AOI21X1 U2384 ( .A(n2156), .B(n2158), .C(n1698), .Y(n1842) );
  INVX1 U2385 ( .A(n1315), .Y(n1698) );
  NAND3X1 U2386 ( .A(n1987), .B(n1678), .C(n1447), .Y(n1315) );
  NOR2X1 U2387 ( .A(n2439), .B(state[1]), .Y(n1447) );
  NAND3X1 U2388 ( .A(state[2]), .B(n2467), .C(n2475), .Y(n2439) );
  INVX1 U2389 ( .A(n2264), .Y(n2158) );
  NAND2X1 U2390 ( .A(n2235), .B(n2057), .Y(n2264) );
  INVX1 U2391 ( .A(n2120), .Y(n2057) );
  NOR2X1 U2392 ( .A(n1451), .B(n1799), .Y(n2156) );
  INVX1 U2393 ( .A(n1629), .Y(n1799) );
  NOR2X1 U2394 ( .A(n2407), .B(n2445), .Y(n1629) );
  NAND3X1 U2395 ( .A(n2225), .B(n2061), .C(n1258), .Y(n1451) );
  NAND3X1 U2396 ( .A(n1964), .B(n1601), .C(n1705), .Y(n1681) );
  NOR2X1 U2397 ( .A(n2395), .B(state[1]), .Y(n1964) );
  NAND3X1 U2398 ( .A(state[3]), .B(state[2]), .C(n2475), .Y(n2395) );
  NAND3X1 U2399 ( .A(n1679), .B(n1601), .C(n2218), .Y(n2353) );
  AND2X1 U2400 ( .A(n2305), .B(n2112), .Y(n1679) );
  NAND2X1 U2401 ( .A(n1685), .B(n1299), .Y(n1974) );
  NAND3X1 U2402 ( .A(n2072), .B(n2116), .C(n2476), .Y(n1299) );
  NOR2X1 U2403 ( .A(n2471), .B(n2159), .Y(n2476) );
  NAND3X1 U2404 ( .A(n2477), .B(n2478), .C(n2479), .Y(n2471) );
  NOR2X1 U2405 ( .A(n2339), .B(n2407), .Y(n2479) );
  NAND3X1 U2406 ( .A(n2463), .B(n2464), .C(next_byte[0]), .Y(n2407) );
  NOR2X1 U2407 ( .A(next_byte[6]), .B(next_byte[4]), .Y(n2477) );
  NOR2X1 U2408 ( .A(n1807), .B(state[1]), .Y(n2072) );
  NAND3X1 U2409 ( .A(n2155), .B(n1633), .C(n2118), .Y(n1685) );
  NOR2X1 U2410 ( .A(n2351), .B(n2445), .Y(n2118) );
  AND2X1 U2411 ( .A(n1704), .B(n2235), .Y(n2155) );
  INVX1 U2412 ( .A(n2159), .Y(n1704) );
  NAND3X1 U2413 ( .A(state[7]), .B(n2467), .C(state[5]), .Y(n2159) );
  INVX1 U2414 ( .A(n1832), .Y(n1675) );
  NAND3X1 U2415 ( .A(n1847), .B(n2214), .C(n2218), .Y(n1832) );
  NOR2X1 U2416 ( .A(n2446), .B(n2411), .Y(n2218) );
  INVX1 U2417 ( .A(n2428), .Y(n2214) );
  NAND3X1 U2418 ( .A(state[3]), .B(n2116), .C(n2475), .Y(n2428) );
  AOI21X1 U2419 ( .A(n1455), .B(n2480), .C(n2216), .Y(n1669) );
  INVX1 U2420 ( .A(n1293), .Y(n2216) );
  NAND3X1 U2421 ( .A(n2305), .B(n1250), .C(n2056), .Y(n1293) );
  NOR2X1 U2422 ( .A(n2416), .B(n2116), .Y(n2056) );
  INVX1 U2423 ( .A(n1847), .Y(n2416) );
  NOR2X1 U2424 ( .A(n1476), .B(n1807), .Y(n1847) );
  NAND3X1 U2425 ( .A(n1258), .B(n2061), .C(state[4]), .Y(n1807) );
  AND2X1 U2426 ( .A(n1982), .B(n2085), .Y(n2480) );
  NOR2X1 U2427 ( .A(n2361), .B(n2445), .Y(n2085) );
  NAND3X1 U2428 ( .A(next_byte[0]), .B(n2463), .C(next_byte[2]), .Y(n2361) );
  INVX1 U2429 ( .A(next_byte[1]), .Y(n2463) );
  NOR2X1 U2430 ( .A(n2360), .B(state[1]), .Y(n1455) );
  NAND3X1 U2431 ( .A(n2116), .B(n2467), .C(n2475), .Y(n2360) );
  NOR2X1 U2432 ( .A(state[7]), .B(state[5]), .Y(n2475) );
  NAND2X1 U2433 ( .A(n1493), .B(n1495), .Y(n1276) );
  NAND3X1 U2434 ( .A(n1938), .B(n1601), .C(n1705), .Y(n1495) );
  NOR2X1 U2435 ( .A(n2446), .B(n2342), .Y(n1705) );
  NAND3X1 U2436 ( .A(next_byte[0]), .B(n2464), .C(next_byte[1]), .Y(n2446) );
  NAND3X1 U2437 ( .A(state[4]), .B(n1258), .C(state[6]), .Y(n2406) );
  AND2X1 U2438 ( .A(n2235), .B(n1929), .Y(n1938) );
  INVX1 U2439 ( .A(n2104), .Y(n1929) );
  NAND3X1 U2440 ( .A(state[3]), .B(n2481), .C(state[5]), .Y(n2104) );
  NOR2X1 U2441 ( .A(n2116), .B(state[1]), .Y(n2235) );
  NAND3X1 U2442 ( .A(n1945), .B(n1678), .C(n2272), .Y(n1493) );
  NOR2X1 U2443 ( .A(n2351), .B(n2411), .Y(n2272) );
  NAND3X1 U2444 ( .A(n2413), .B(n2350), .C(next_byte[3]), .Y(n2411) );
  NAND3X1 U2445 ( .A(state[4]), .B(state[0]), .C(state[6]), .Y(n1254) );
  INVX1 U2446 ( .A(n2278), .Y(n1945) );
  NAND2X1 U2447 ( .A(n2305), .B(n1814), .Y(n2278) );
  NOR2X1 U2448 ( .A(n1476), .B(state[2]), .Y(n1814) );
  AND2X1 U2449 ( .A(n2474), .B(n2467), .Y(n2305) );
  NAND2X1 U2450 ( .A(n1946), .B(n2240), .Y(n1961) );
  NAND3X1 U2451 ( .A(n1982), .B(n2022), .C(n2204), .Y(n2240) );
  AND2X1 U2452 ( .A(n2066), .B(n2112), .Y(n2204) );
  AND2X1 U2453 ( .A(state[3]), .B(n2474), .Y(n2066) );
  NOR2X1 U2454 ( .A(n2481), .B(state[5]), .Y(n2474) );
  INVX1 U2455 ( .A(n1751), .Y(n2022) );
  NAND3X1 U2456 ( .A(n2469), .B(n1456), .C(next_byte[1]), .Y(n1751) );
  INVX1 U2457 ( .A(n2445), .Y(n1456) );
  NAND3X1 U2458 ( .A(n2478), .B(n2350), .C(n2413), .Y(n2445) );
  INVX1 U2459 ( .A(next_byte[3]), .Y(n2478) );
  NOR2X1 U2460 ( .A(n2464), .B(next_byte[0]), .Y(n2469) );
  NAND3X1 U2461 ( .A(n1258), .B(n2225), .C(state[6]), .Y(n1800) );
  INVX1 U2462 ( .A(state[0]), .Y(n1258) );
  NAND3X1 U2463 ( .A(n2227), .B(n2069), .C(n1987), .Y(n1946) );
  NOR2X1 U2464 ( .A(n2342), .B(n1790), .Y(n1987) );
  NAND3X1 U2465 ( .A(n2465), .B(n2464), .C(next_byte[1]), .Y(n1790) );
  INVX1 U2466 ( .A(next_byte[2]), .Y(n2464) );
  INVX1 U2467 ( .A(next_byte[0]), .Y(n2465) );
  NAND2X1 U2468 ( .A(n2340), .B(n2413), .Y(n2342) );
  NOR2X1 U2469 ( .A(n2473), .B(n2339), .Y(n2413) );
  INVX1 U2470 ( .A(next_byte[6]), .Y(n2473) );
  NOR2X1 U2471 ( .A(n2350), .B(next_byte[3]), .Y(n2340) );
  NOR2X1 U2472 ( .A(n2433), .B(state[1]), .Y(n2069) );
  NAND3X1 U2473 ( .A(state[0]), .B(n2061), .C(state[4]), .Y(n2433) );
  NOR2X1 U2474 ( .A(n2237), .B(state[2]), .Y(n2227) );
  NAND3X1 U2475 ( .A(state[3]), .B(state[7]), .C(state[5]), .Y(n2237) );
  NAND2X1 U2476 ( .A(n1993), .B(n1963), .Y(n1654) );
  NOR3X1 U2477 ( .A(n2351), .B(n2350), .C(n2461), .Y(n2062) );
  NAND3X1 U2478 ( .A(next_byte[6]), .B(n2339), .C(next_byte[3]), .Y(n2461) );
  INVX1 U2479 ( .A(next_byte[5]), .Y(n2339) );
  INVX1 U2480 ( .A(next_byte[4]), .Y(n2350) );
  NAND3X1 U2481 ( .A(next_byte[2]), .B(next_byte[0]), .C(next_byte[1]), .Y(
        n2351) );
  NAND3X1 U2482 ( .A(n2225), .B(n2061), .C(state[0]), .Y(n1637) );
  INVX1 U2483 ( .A(state[6]), .Y(n2061) );
  INVX1 U2484 ( .A(state[4]), .Y(n2225) );
  NOR2X1 U2485 ( .A(n2256), .B(n2120), .Y(n1993) );
  NAND3X1 U2486 ( .A(n2467), .B(n2481), .C(state[5]), .Y(n2120) );
  INVX1 U2487 ( .A(state[7]), .Y(n2481) );
  INVX1 U2488 ( .A(state[3]), .Y(n2467) );
  INVX1 U2489 ( .A(n2112), .Y(n2256) );
  NOR2X1 U2490 ( .A(n1476), .B(n2116), .Y(n2112) );
  INVX1 U2491 ( .A(state[2]), .Y(n2116) );
  INVX1 U2492 ( .A(state[1]), .Y(n1476) );
endmodule

